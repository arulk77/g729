`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN4jZ7PX8JDRIp6s61QCFzCiHogDCwGdti/4thAuhvHVa
9uVCUQmN46+kjgYkyizLtMppd02oGp6jzjtkNzlJ17S01FfqHfWGU/Ye4q5am5Pe
+H1WGFXmKG+q2LX7aqWNtwMS/U+CMrbeFIuPp3dFcimDeimJy0w3aeeqSeLMC3sI
Z07QYsWWizKAWO57Qasc5GyEiFGpdVPyrh7wLAv2+cu2Mgl/YHlssh8D2ntuu2mP
cKwl/XE1+89QTW+JCqDh9verRjQxFfO2MN1muceXOptTA8u/FXGEF1M7ZSRU6RUX
eDSn7ZILGYhEhvRKtR+YipL+EuWYDAh7mxoOexlAxR6ljoBoPovxHsYwkscJJRYu
Zx8ZoNfR1I0S9gXd/a+AxIwuMqZolcFJ/023rOcMYx3qNWNFLlG/tGOq+IBVKUWN
6tiKi5hhEZIOL+XlbfmztqL1wkoG25MM3IrPwpjF7b/Szm3VZFYko2OBqHeIVOT+
Tk91gLqk1C+33nuhY61811lDlho407nLlexDjmQFueJBM6ADd4/R4wlahC7ZPqxT
/o4bTwYZoM+P9YRDGIAomOej2qfFifZau/cn+PVrMTaT5KrJxIwyZT3EnT5z1sXo
jjCyzpiY+tlR1/8vaN1/Ah3Lbz2gGqgl3iQl01zP75wzR+kHLEEHYq5zev6O4FTM
GR8G/3FMe0cGyM6bePcnBMTO9xSaHgASwRjzM+zoSiXxJtV6Cy/WZn2HbKYa4l41
+2pxValwZzUEVdqJ2FNCweqiYzqywMNXBg65uTaG+bR5FcYqEjpgm3b2/WhTyNbR
xxJy9nVWXkao2hggCkHlTcuBEf5rFq1k1raXE6yhv4zK38CE+zNtpKQ3y1+ZCph2
H1Ko8DH24U2ZE0/yduM+ZZX0aL6TrqnCGNY43rcjq4qs90qQGK0vgeLGAWN5tz4Q
uh0cSuWLV0W1W2/6QIF7nqabnv1oTRzSv0vmVETCUSY9BS7RbUYaEIrgJ9mwtCk+
2FdKgkkKP05TlscjlYQrsM+bnUwxyq+7oICBUI/n5MYB73kquAPHAgl6VI79X95X
9aPLXldymBdCHRud7bMA75wpgGKHKH1NbvRz8fsZDveeRSsAWoX2ZkpvxHPMgGEM
WOoJM5ZJVw2fydbMpIn91DnKKF5h5IUdaxYGEaq7Wajy6F2oGQ7BNnKOHp+JSl/a
Xir2RpOnL+GPffvmolTi2NcDZCwSepMqv+dfAzVjYjHyPOpeoSGMsg7Hf33mrSEO
yM0x6bgiK8TVseDWULF/kI2R9piLd4Ns3PpwUX7mOwpX/qNxkkqrBGjnpJNz6exg
l74fX8fZwLhsMLbVIldgaHdCgtVcJK7vSKPVVqjDnkU96OzvjEdRA3a1CUx3V+um
U5A7RFxgUZyEGx+F6w6ZQ3IATxc+EC54rVq3A+4hKmZWwVOyskhSYQxGkEvpr2SY
JAwv2pr8z3Osmn+sl2N7hYxHjxAiT9fi0pxyC04FLeIz7f7bc7FcUswvBndq3voN
UZL79zBisEp/mbm0UBmzoP6YAAMqVJJT+lkiqJpw0M0LBgKAf3TC2k1HSOVuhkji
WXu8ojhKsAtS5BsUnVRFYwKWnuV96REJttKZ0UFq6CZ1SCzlXUCEXlRZDL8TLX61
bndrbDGifu4msSxvx33DTpjTa+GX2co8TghCt/Im857bJfMZS+3QNDbQXuoZUnt0
FDURGnxOpACcs6z3sNYjVKWBUdZYtQA5pjFD71Ypb4gyBlur56eQABJcGeDAC48K
RcFTewkf1WeksXVPtBUpZQILdMkecuE3yqUCBuM5oZ/5ya81sCpuu4qEQIcFR78b
u8h2VmmEZ97tHilbyEAwkjYfYjlNb/79/SpAhuirs8JT5WpskgyiFK+1hagTzqI6
Z5MG8etGWO2xCN9AOTklQoG7TuRKCOgzZXC/CON0oB93Nv3ktyJLqKD++GU49BHF
Wg+ahGfBDnFb3AvIOmdN6fQIvOpIBJZw/pU4Q/k5W9LYSfIPm+G1BgbnsXj2+34v
EwTwem3cduBZoej/E6e8mWBzFBBdf9uhaBmcWzBwkLISKI5j+tbM38cK1M7fjAaZ
nf5OMEmQzTuGaQjY0QVFtq+S0W+wlgVLR4hNkdT5oDr8qNbHqqWPv8vYTbIxXSRt
H0vvBkX1Pd1Mlca00amDdnXMkLGsQzdNVeAWPppr7BB9wNTKzd9w3IusU4PaB+ct
uZahOhNwiqLSVn8wjsMGnwS5x91oOuKajbFSKjeSuuQLdQjYXj+1tZjwRyegP6sX
zNaK9nXcw2uiGItMC8PRy7375/TgE97bFxbbz/n245otrrMmuM8DZT1xD44lrrvw
YLiC4LesCqSd4MXjFreVcBmY0FkfX4gwTaBbuRS64lRrFbBG7u2qVV80EUp6W76S
EVGPv0QlIm5SphZZF+OOBpm141aEV3HA9XNdeEiVOUKK0j9NbB/owHA7XzAVlrpF
aPBprHhr0uBj0OKhy80lXLy6BWGGAmdOj9tOCa9tpHmy9wS8gajCKqBfjqiLnveW
6I+miYiFRecxjlKtbfiKYSMZ/Nf6Dyc91ugGZxSpMdnt+Cs2cEINXnUY8F9wsXld
kRvqtVTwEGpTrFJYaXUlcxmhLoMXcmUK1qbBb3OH6NRXi8HAtg9agSVc/z1C3r4j
ERerqkEG6cpKqFKLr+ZDWu+2NSoOf8liK9+Yi8lsRlXocZl9vsXjXdE3g3niz5Uc
kLxBEPRaG6u/NWiltmpbWCRdyIyfC0uXTjUyLbvESw8kvprZquP5ZdxB891y8BO9
5s6YNuQvRVixE5lHUMBe6K+gH/m9iFRx2YGHsMNlAauldxBtTTDFQD1Umx75tpRy
fu+v1iDPzX+x/teMf+QQSS2VtcXbxLACa2dERkb1aN7qPW8EnL3d0ZNt4Q38gMrF
n3qpncUlrB6RqBq6pGA8oxx4FenSpaKvRgbJK7YNYYVIct8s1PgubGtSmUbCBgiQ
7Dc6agsue7ZGqGcbThiEAncLXT8qaZVPFDylDYkLRHmtjPVBCDq4liRiXNUXqo9l
6/57lJ9kJTin/pjo2pO/0qVOjfLt6+7WFDsNlyNfDx5Nc4tMPvcK0NIze3j9Hboc
MEtprjxh3QA+IqHbFki422DI57+tBDNZ6Ikl5T+HJhDzEzdHUCaUbNGmJx+DimHG
k7JakEKcCcQ4r8T49Rxya/bqZjjVHSaHp0S0l547qY4/DQCwhfZ5j5+9W9krcM59
23M/3hsIjBpFFP9mc5F6F4pLyL7guu08BzBBHtWRAka0whWuOo9D61RmHyLX5tka
Km69pzuXlL/+j4zoLaYxFA7XSLGDE/+3jyBEmIze9f3FfGcjahrJt/wD0LjOYeQS
jM5PKusbDTJG3mU6C0+EkdQ9Io73K5Rl1DV0s4KbD8dX5CIB3VYkrip1Z0h6KauQ
gQmkHRApSZ/f8GVopWMkTyh1tg3Kjy8POpaJC9Ekd1SRESUFNruPQcZrpXNGzzwI
y7zSvJdvDBeSrdrcYe4RPTsbflr5W7n2gRP1uKwI3q+S7XgEpZAONCK8EJ2/hZqI
g60RQVaO7Yu0NqQYcLNtq3xLvPCErit+Bjr35b7/4/CfuaX+K5ykmdNS32nU+E7n
X4Zo0/DuYR+hf46z2qvHN3Nu31r5yVxR86GlFssGsSxNHWaa9YSt02+dCPVJTrhm
E9MuJlzK4cj+OS67j0Iedts7UTZtgcpy0QDUFy9G/PrS4sUgt85/Vsb5sFYTLFIk
FM7W+lh6iVoVTIXIAeEfntNH3Vj4cg06pNH/yMieKsSTMyn1ExOcv4zxw7T7/oGI
gu9EI8VqmvX4fOvR0RsoC9Dk4CLgFA+XwFXa/ZvOKl7N5PyGEU2Uqz+O6qGRUaRO
AwzLlOweN+ZLPAgSnMfs1E6SRtXBSsS9OYgzwaPZbV/Q/DXSVhQCUQPZ9dSsXpG2
cCD/Zv3iThCmzNjxp+Gf8jwxFT2uWmaZBMeajcjjkxTiAPlIN7EiVbIzgoJ+DtOB
Gr7uroQ/yXfFfqjtw6pWtIIZ+aeptiR5ELJ9Ty3mJNxUi0cgO3VtURvWoxXoEPSm
KOXxp1rU8hjYoJ4epzwoCY8WG4DJz6DVIY1lg1ku8DSvP4bszHxDYgRIaOpfsZXA
LJKm1Izp8r8RM2SYcskB1nGpudzUTrud4gqnq2s+6JOkXUBoMLp3g6dVprcR4kgA
tIbfriIKTX4WznL8hUTf6Jo9uZYP8fgQ1iEmioKQkHg/GMHS/rGjVNgEXQbzFkS9
AEKRfykUsvewDaf3wq7mCDGCGgZ8++up4xsS93Ey1wGCq54jLabWtqPD2MfYEIGN
elAWZwJF+pcr9WSLbMY7LkRukoyayqwsevNH2boQnVCX+ZGXlqVY7lqxIsP5ifOf
o8smy++GaoHvxV33j2TBhwdtIrS0CDqc7gqKJDAxA5sfOIuI9o5ASX50gMlVlm6x
LPEOJqhBgeOEqOBIgRpsFJuJrCzzpIyGsHsaUGbOjx8f+vUGdfE4nJbRYeOBHVhN
m0qaEEtRQCZqHwNMy4AOMEd+aAlakSJmGFgsGXx4XByfyrbqXzS2Jd2nRpq2WmQJ
ay4sgpkXRcjmukC1zGEgatrQ1SodXP82cSCuE8TrBinLL4zvEmEtCAD5swNh7EM4
8qt5lBxFPMYr6wk1bPag+DQQhc4GyiLrBKDQvbEd0WuKl4KHyzME1Nm1/yXAGaT5
GEHoBeP/0Nl1diaz5mLrbtGe3uocOdIvA5eon2W2pQekTBDiuka/8jfaHffYio0b
2itbJBIu2ydPBrieJn0B/QfxS7m1i9ALuDXBmHDJF7MSxpDSVMwMQjkUO/EXLmza
8HeSO5VCFWMzTuFhppku9pt3IbugCAymZRNnEzigs6QyTuO1uoYJjwW3gD1BY6aO
qrfcjP3pqHcal7Nu4XMmN/TMQVAQb86faOWz595obktFU8g+WDHwE1Lpo1/AcJVt
S02wIA1DpOq7xFz3if325EKHHVihuwOrDfMA2tVR1t9DAbaqbKZa+A2BVfkjnO9i
ed+ScnurAT463qNAvl/alas54piChxAJw8ser4X5EAcjVji+4tra8/5+OwW1cAtw
OTbNO8ptAMfQOFjfiQutIw==
`protect END_PROTECTED
