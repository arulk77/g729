`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/UKI5Q4HJ41IKgkPjhd2UCbpGQ5eSoBlKJ9sT9c7CQnw
6D0f+k6Qrlj3/ej4empeHPKBLhesVnepwsEDOJdUf2FEko3DG/AjK8NwdZsrs+1d
XDE6F8+GVU6dsqWUtUlU/rObRfvzlaSf51JT+oHFNWq2KVjj7xztzvMOUm2IMXc9
oIgylr2XHpUo6D96c2dLtlXjQCHbKyHZIwI1wktHqBoBOxPcYZI2NLkkkeyZem1D
5OS9ZQYEhcHyFMX4ETfEDJluDehhE74cWJ4h1C3z4qNc2ggP6iZRhWHXzjkwtJru
UCjO6JK08zEoKn7XrLwKOPl/q9gIXU7R23es/oBoU2q7aShbxZDLtzSVOmTtvEFb
c7dE8LdCfXiqrC+AikF64PBDSpwTgVfppBJiqHog2UxaQlyL+g1W6KBN8A6FqgZZ
b2Zz4rKoZhVrNwlRE+oravhBGBuR9qSHlJMscy1QqEviR0VEN5o+LJM798vPuXuC
iOrWzZ+LMI5QaUwQEUo6PMluv+A0xI7Ok0mdi0EiAlb6FnZKlAnrGwjzUU0rFJyf
x9dD2mfTsfCtqMmCf31tUA==
`protect END_PROTECTED
