`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44w2KqOkm/su3DFP9LNJE49qGzGLAOUrqeRw2TrlI5N4
1zEd62sBQVcanVfB3ndVoc3y8aFtbUSvhVCS69M+YpzJGgoXDQ3NtFF8uGXdRTTd
7Wc2k6WTb7gddElALYjleutcJCB5a0iQj1w41uBsh3KpSD5MyzmOekx4sD+cD40r
59muP9Pz7BpVNKPJyXm5eFGtpYN14YEpf45MYP9xxhxCjC4I1sSqHp5oKRFXKUHP
Wp2t2w/XDJ8wMqcV3I4+3eVbh14c1N89BCmRHcXa9U2FF5qS37f+eEPCdcQqmB6m
p3ZgiAT+AZioBIscrQOB+miV8I1AUkIwCq/v0pWuijXS1zE69L3U/9RtUvanADQC
N3aDo0/N54lj99tPCkO9wg==
`protect END_PROTECTED
