`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHbQWhwCpBp8e2XLerGqYL2DTE9sgB9lNLA2E6/81ZDl
mjnOAGqc2FKPlYeTEjEBovGJTQUzioCez9cOW230PUxhxY3q5MWvfTP/3dD4s/QS
8fZKfuLJDcIsEcDklqGmx1NjV4r+ivoe5AGyiZ6UzHCZmNLWMiPvF7HhJf4QOrJs
puVt2PDBEloDP+5cnd9AJA==
`protect END_PROTECTED
