`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZBVpOwGlnrSMAcmZ1K90CE2NtqI+r/Iteq/Tpd3gWLd
qm641jp08iSEpbwKJZjhRtvVRrpXtA1J/XQWonQPP+OQMzb8H8aNAgik2bfp4KMj
9m0UjShMpcsa5hZCuOyaKXoC0Kkl+pno+yhQ6BvRBGGcnRFumXe2A0CDu61V+fJw
0vAnq3iFeprXVYE0di3RJyEirPBO41B4PuA6rJMUcaVc6xZVavRbnQLrXD3t2ezX
DTBd7u7bq4Mh+UEOnB0EamX28yQQz3+dQWbzjAjs4IZxjiZ4GG8wVl2FnInC2QKJ
Uj7JIJhTQn7ud2i45WwRpD7ZLFf2sBd8uuOqf8cdE5MOEBIdHf5wFE4ChomJCBxJ
0a8Q42GRA0dqN2HTs0ysGEAejVh0WuD4I4e7O8ZrV/8=
`protect END_PROTECTED
