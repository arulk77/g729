`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42BB+uf5WXGGdh2rtPfpwKdiu5TZ7iLd1bUpZ7u8+Q/A
N7YVLrO0+/jrdQtFqGNLx7lMKkxpsfXeu0pTxrSd0O2/PzieDAhZWyTXzSALSRul
FmKDLYmQhpsHlrUkVvdCna+XKkA4Sv6vklvsVwW9XFzsvwc1ZGoAukXNahMLC3+x
euQ5WN7z41SZFO1wJpgblAClUHwhOQo3i98Rw63hXVIPTFEukkQBDLPDpW5r6jz2
Vcs38LNW0t0Nx+2uOadgsRxNJvlj+cLluQKpf4ZPoRrlKkJonuETHJ6W8AdOvC32
3GvosNl1xBDJ1vpHEf4Nc+9Rb6t7k9epJcseMKgjYk+SvauMUyxtS1a53SHLyyO8
u5T4i8LCNuMuuVGl6L/z1Q==
`protect END_PROTECTED
