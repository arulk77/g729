`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47E+kh0TZN9TdAxS6XC9GICsC4ZFsQV14RbTYWjf/ye2
pZOExLwMNPBzV4RitCiPfBOYJG1TiBPiK4kf0Ouw1WfI0nu5ezRoIemkV9XLmGCJ
WBW9sBKY0B+Vo9t3+yPpasKtu4cs57/ORvzwkHKRxWQ2WgsIL1WyqhnYBVMI+BPW
ZqsjfubDIfsIG4RGEYpD2ywJNSekclYna7w4TuP2FPU=
`protect END_PROTECTED
