`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB5r7zQX6z0hvRG295kfZs7pbKrcN0p41wJid01FvnVh
10aRvHDQkt7Vq8KjuWfmapJQZsWOvNP0Wb3eyFnpMspBwE1zTnCyluucWgq1+Wdv
vZzJMuZ385xfNAbRQ8OtFAumO3utSKt7mwGxoiEJerMFZZ3E78xGf4MzAzngzj2D
GPhxqjZ6byDJKYyzY5Ga4CM68+oYMLRxiCnwGHXlFDcrXWKlvmC+PiS0kB9QJ9XH
vmJcqLnOjzUBtXFs6UoI2aGi8pAhKUTpBpjdSnroyuOEX8IzFZVAVXvDN4P5LoZa
BVOHYjch+SUMDE5rt0pKcyRgDqu20TE7ly7btnquNg5w5lBz1DkcmpJW/IV2LD1W
eDA3CrP8hkSzrwLNmwgBi5XJ2ZBiSAD5sGLqEU/ijxZ2Ux22sH52CWBXDVPWFGmi
KjPmO6FpJ6OgOvjIT3EOSkUVU+eXMVQici/vhR7/F9rcCvoXHtwoqnto5DzUcpwO
6OCH4jCXUC4TKfWAZMoWftfSjMTdoz8r+CZgRhxBf5LrfFjSfqiNfiO/ZfVMhKCX
9B+HcF8EveaKvYG+bW7PON9unK9ARgaiTaGVfR9lVU6q75MMqRUO5+deVfA8chp8
GG1UcCIvn7lU9mU2VxEMZFzVPfp0Lyet+HsonvCZPEkc25auSaGUvIeVF3M7vDEj
`protect END_PROTECTED
