`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOyrPdOnCIt8JAMf2ZN+sX2MWcfQywKmdYop9yrRk5zk
+V8970QUX4W2DQUHZ9+PJQSUoRKiXLbgLLw+4q7eIUhVoyCnYS7F2KAm7KH5LnIW
jzHcb6M3I2JTpVB5/eObFKS48OSa4U5anq2cF5H/KimkVyMOjFIyOrC4kfO7JVza
Yho79HdBp3IeXoN44ItQ0inB7ue6c7zo/As0ImTlSHGUpfidd3qmv6t1dvPuveKL
Jpk7+vvw+PG/m9YZTUDH/LzbL3LofJJcmun1NrlGTkJTkzzjTGWOUkTqcbkz9ofI
5PM9XQVSn2ZgMSMLHA16Ykc3J+KHgwyuWO/JYiCHObOIyBvQaCZb49Omtc76kjiF
uQEpUNBZhhHBWmJIUFCuvUSB4Fk4UDMSDCQp+pYoZ98Wc3GZWTE2Jw0n1K+CsQcP
c+JiInmO5Ys70edM0x7NJG2rhD1nPQ43XjbodpFm21XhfIDWVHKOPtrrYNAI4nTs
`protect END_PROTECTED
