`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHprz69LHVXp6hM/iYDrqp0tU64bixacTD/cgG5N71XB
04vCM03A+OPveb8CWP/AMMpnWXmO+BiN42i8GY2+m48KhyQdbiiXv5xIRUkF6By9
lyjMWSV58/utJSm7wPWUsONEZkT1NXnWL4q8xdKyDwN1MBMfYHfsItkL60PlXL3B
AGbAZ/c/UChe3W9KXg8+YDTI9qDdpN1tmDr6G00DHSPEdBKS+HY3Hq+3VrlNDrJ0
6ape/fltRcEFgGSIq9PdeajNqQaq5CxrCiEA2Wd1L8UetfdX8hFKEm4xPjnshY3o
R/cTu0Azrya4IIfVRiG+6Flrd0EmbGuY237++5Dr8hij+WKnW3Vo3ASxDqkgG9DZ
`protect END_PROTECTED
