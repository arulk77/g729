`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIgCcZic3dfTPOrVxPzEbeXiNCsmrJpDy7qQmr43AaPO
kM5Xt4N13ZUi0avx/IWbq75yyWn92gW9vnvvFYeavwISLZtxW7z1ns8s+lxBfnpq
y7tsJT6yECjZk8B1WX5c6NToxiGZC0lwgqxDV0X3EwXDIYydIHGZdzXQUxhELovA
9jsKtRojIB7Fciixwo3NAtMPAjokYyeHisdrYwsYJbSrt8yW5DF5TG60vS1w2hZ+
uZuV8SetSEgS1cIYwzdGjz5uOZ2+Q68Py5PF5GkXAezbkw1t8czHNR3fEwspO/Xd
4radAk4bX35P7M6WK/j1qSCNfklUTuCSbkVXExrsU5mWoK1kMgJ5wMafkqtIKu3O
`protect END_PROTECTED
