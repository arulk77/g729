`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKYj7W2p1m3GuQMWInR8Ts2be53cVWLJdWI9D4owQrUG
eeISecz2toIZu4yDSSdMeWyQEsUjNS3zPwlKQNR4pJGK/lYPOCPX5MMV9KTgKOcZ
xdNoW3tSV9Weyfr1HtGuOa1951RKhZ25BTUt5k5a90psr/Vhv1lhFq3VpoeuVrGj
ZiNKVU/cVhPLtLQc5p9/JwQ8xFUJhay1m66jgEvFmQQh8Ix/JssiuMqxtbbkO/2I
`protect END_PROTECTED
