`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOwmlrdmji4xVHDXhCApuvbAWQM3v6wd761WILv3gw/n
nVgYLJnDo21f9IWCttDaHc8nKHPwheFO/a2QTpFCy5oxBCb54eq0r8Ndis4CpqLF
KCJqD3kjLwvOK4j1RKt0a2YXyJYdyQColUOQ8sU4m/fvwUbjKQonT+YD5T+G0cdE
QlxQ1Sm3grzye/BnzseeRNwUtqHHa1oZWT0phDNVjVJf7500ahA4GZcT1QmBPlzt
`protect END_PROTECTED
