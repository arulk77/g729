`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGrR/yYLebWAq0j1Xt5vXa252yTR5E//ng3IHVlXnCtD
YXw3+INr48WSnrjATh84j5UpPxPahqmMHsSZgLD/Y6VzlUTFkz1e5JBeL27qm7Ds
DfbuJHcNa8E3cAqsqHQODuj19bpI/DqUlC1EljwewUVwIGOfrEXnDoRvCp8aByYe
m4DRbqCmfNBOWLwnl9H/vpkzYVIcbCQfd82d0jMh88GD3D4SuDbpRBCTVC6/2FHo
WMZCizCBG2O3YuZyAP/uAftMa00Wj6daScckD3tPvj2WxSAx0qv8xxBv47niVFfz
YJYDKu42ezEuo0wFeAB6Vo1ybPfI/yx9iXzCdLvtZChktUbrQX6M/EatncK42Z63
nE5p8VuvuqjP+R1Jrl4CSS0N4sv4inD0L/IWtqW03R3vVDrgCiKgojCMMBjoW7w/
lMVYkxw8Jg8YDE/afFIxFfx2NRa8FKkMqOvQkBtSe0k=
`protect END_PROTECTED
