`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG7C6o54c1WJNbPEac47Dz2BKzjY1eM3z5b/wzSGrtD4
hIeaGJ8uItiy+Tqd3+i5syqk1Ligpah6g/s4je0yx0NWbSc2WIbkiVMjJo7p1A1/
y0MOj0L07h/jUBWAncNtuP3spQFPYLvM5ksyT5aPALW8Xy3IAl7yhwGYsJI73+0S
ZE6J/1YVpKINNIzex2JCwcdWe8XnGbVYJ4tNIej6X39V/FJGi0aBHn6NjvmFZRci
iyceZfbib8U3I6qIjKao3qduHrBL5JzPereCnytoN3HCNZhOgTZV2FxxkldJRbNm
oZx5HRS0f16b4BG1R4FmWuOXb/G+rt3ap6wOCczkFnVa7i/2CVCYvGpP5OiLQXhE
OmYtAcnIjyps0rE1MTvYfhvANSgzaYd7lW1zLTV0jHcJtHWQg5Sgivnfi91MIZpi
R6fR10BLKJfF1JY9DkikjqKztSWQe5Xi66snXi3rAhVAU5pIAv9ES4lgLZVANEhK
`protect END_PROTECTED
