`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
b/P+zNh3zESg25UqazXzLv4N4vxVzFntrdNARzIAB9uW5AzJJawAwws2A2vSIoni
r4bNk5z1hIt9zAE4fCmWqkibajJ+8Cs27uE8n6owh7kEN7bRj3kX1+SS8C/4bMDR
mC4ollRBAOoVOBKKXqQDtegrzckDydVFY7p17dNnclc2k30CRCBKAtOq1vtQ+SJh
cU+t+cNg883bfu5ot4qoM1xQnukSwNvOwHL3zBBrsLK4yor6j2ta+JotJ5QWGIbh
DJ7KY/+OILQ0M6rlmbNBvKXr0+x33GCcQkbzGTx0q460JYyXVxXydY0KBmQvczzo
tS/6wlWUfdrKXze/ffxXBq6KERDgnLQEPZTGHkJSSawed2GHDm3UXDxfRJwUCjzH
Qv1SM6BHCmhKRa69W9+wMeiqaGrP922vp4a1wei6eh6orl3TIRgiOdAcuVI83bSO
mg6IYxKITLLIJqdS4jIRV4BIYzxg9vAxRzIbouZSUyIW4WDiwkpR2opbybCmnrbp
A/AM+sdZP0x0pce0wtbCT5GJFvoCzZy9U+NnWh+R08CiE6KUeTVyX6JUnXJGG19F
ZDi+jIVE2u7ERLwyLBaejNsHBlBGWF+H+rCBDPQhdKqKtTx7W+14EK3ZiSvwoK/E
I/Pq7tdOP8/L3E+IO69HpJppn3QYXTBim4KE0NmYZW73OkRutLAHCklYnBa16UQ2
DoWuMzgDYI8CQJQ/zXF3IkD1nC2NY+XzQyaky0K7mZBOLzc6qQ/M8d4N5Qw1FFxW
FjH1xbyMGgwkMXM4Gp4xAdL/GrawkzAVZweRs7P2TSFCZor9JxNs4HI2lOmcpVza
o7i8rB0dFXP8t3fg6uT67gAUcoXYoBf+eWDVzjyu5U14LZ8Mcd4tY3fjfN/aanIJ
Eh+oIwaItvJXSmrhmNelQe17kSIiU5VBuIn17rfaU/KGqrh4k8/NZuDXNecSWR4z
w3XTKA0PO85ZaaMPesG64bNq8/XxF4EkK+ubr3nImBYUZYGve2sk+96PaPVjkZvd
gzfvSFcGKycE1gQXPnGhHm0XuYGKWwhLuoSLefW7qzS5mpW2SmTWL71whfiFJbut
gZH3klW46tJ3d8sOj6d9GeM7JlnVBDnB6WY20onlxbyF9O3MF74LGrB+hGKrF+OQ
JiqlHlDODQ0uoCipypDt6HS/vAArzYZ+R5TKEIiNT3+3a+CmO5WxYn3n2Fr9vitS
fKZr4H9XPbjY1Hjj7mrdKSRjmudhDo1DHCYFcR0n14fYkyKZqT2o+WHAwxJOIGcv
3UNiH8gGtMgQPH7zvsiAKwsIA7kWpLIWrD2hPNSDPcIf4m9/jL49Sjh6YKjTHjhj
IlUroH2AW/URENLygOqMYcxESekEw7LtR+Cn3So5lzdy5lJ1Yeecyu6Iqr3M6HQf
jCzSz0OPr4isHcCt+iq5s3QY39TTFnFaezP1NlIFLi1P0L78f3fFy6iigKLYYZse
nGJFsWv0QSfJkP3gr6b9EDfKs4PDUiAKzKYTlI7YEQ6fLdHqGTthrv4aZbU5bnol
s4TH5dopoomuz9QNwvamdMcplsPagcGo4D81P15NFL0Z+hziModt5a1aDqBPOnCX
iiJRomJB5yNIynDxpO8OHza4pxChuh+j/LzCsXteBayCVrz856YbLVfWmNH2Nr0X
B6pnlTyE9AkjPw4Q2O1ne/d/K9Ma8PP+fGIW/w99iarh/g2KXKGuCk/Jez2Um+3U
rTDNG77w20kZZlnk7Gz1Gvju+XCirT8M40JolfdOCOsAFzFJjQCsmwmdOpkr07Uy
+7xibLQfN9szzRguRu0qk146Y7TtAPzQ7TUZ0R5tacLi/356SPslQGXMU8PsWlHY
lgPB1RNkVl8vkXY6MNnph7+B40cXsT3UvwKij1tZIvS8JkBI66LjZeB9CyslhQFG
MkEewM/qAUyjFQoGiX6isVgn27+G5hZR0r4HjPhzYjLFnaGDEIQ/Yug1IGYmoMeL
AedLtnPaSE5vl4nMJfkJTcT+W8/v7o1DMVMx2ywuqLsfyP14/ax4z+Q99geERL8T
PgO8XhCOuURrZvbadQoFIqpVdJxSI7DgcR0R9ObY1nbKZWo7jA4Wq6cuB7rRcDKn
ap0GQyeMJb8lfA6FLYa3Eg4YJo+wkVpyui4hHEKtgba0NPxQqBM0TtnVRidTOwB/
nQgIKGHEdvnnPo3PEmbQVwtDPr/O5BB+yz9yZsJ+w03SdyzkkF5Na7ingR66uivD
Q9vqS6qbv9X1qks/Ssos9Rd0aOpVxuysP46rva5RqA15o1s/Ay3OC0tIL1m4gyzf
IvG2AnwasWN4OOJeYaAQ7RL35GhfTOScICD0UOpYidHhq9+q0LVrniVBer0vxLsT
SeGdpYwLq4VRjDEu2nfs5RT+VfAgtChwRXJoJ6i7H/pUH4J5c3I0RKUm4SzaaPSd
vPEgbyMjCZ/jGPWvUvEPWzLckAownaqKvrw8e0x0d04m9bpleltWBG7wHvS63UQy
6GdlzOjVXUf+mHoIUjjCN3SVOONA+oCixexr1dDklIDgFCG4xAdPChKDUuKNL1O2
ASeASuZAC9kxb3AIvLkuiHmct3FHkylHJnUYx1pTgB3vyfeGSyQ0xbuDNjjpRta4
o2Iw9Ks/JjWONFZHM52kYFageYnbCcGq/Zgwyt8pj/QXxGBwH1W4bba5a3SBCSIy
PbAcBFWulTVK5dxywGkaOTfA9qFX38Dk5YOXeiOqhxhWq+c8mSxY24mqadlKvTaG
7hdM0KFlaUwU0HFBrZyMuh5WRGNyRbUcLJ//lyue6U+gxkm+CqLPf1NutnTuhQN/
eagqWB5vUAWNAL5hygI0dtDBR8inFAVC6WCnblolxFW6Ph9DymiPjIs5ewwqiQp3
1LUmdcnWS5KcumKenbX4E3HCXiRsLqViu8SyNyHfMVQzNyT1QigluDCVwZmxTqxU
TOfGIKtelAqhcScxviv0Bw6sHeYJyCoK1buI7OXIc3R2D2u+HTrXv8KrKAhvm/ok
VGPgaMOSCImKepP3DMwZACHbOS8lyCZ+mQGCQVikfxxwujgM7kpYrT+NThivPVce
x6bjl6g0srpAqOIbJiXEKamrcpRjN1XyvNYDzjFGAZrRYvxDHSZ6FITGBun2+dx0
tCRuKzbb/7Ss9UbQUrQDs1UC4xPUGPK2/2k1ZS6msASwDRt/F8xxHaJ/Eg42NSE+
ocgnsJckFptatb3a5fTc5LDitUrKm4/5qfG4FXB9M8FuD6A60UmAcJ7u7nwswq6w
7xsxVRwv6uuC+5piKsXn8CUq66YDdSFH5cFz/qKkVc48mPe3vJ66kZRMmhc8qdaA
p+xPaNP34Ha+7/IBvdK/Cmlo5nUNtM3rPVAL+p9aBcRABYXum1PWbnKKuKUh6k/w
Mbs4KJ703PN+xIxgUOPDR067O5196YugS68fwn9smd4u6H2SBkSP6AJiUb+2X3GM
O/fQ6VS/EgWmc+FYpAuESX51wpT1v8lb6+TIWNpF3HKeExieOKwbvcKZMT+hNPBM
kZcl1ECDJUdxhrBQ4EPLzaCmvOlZn35CpfsZ0lMQktAGsTj3RI25Cz/0pmrX3dxF
xZ/5hkA4QgGW+8wIUuA/VXTdfdtUzUGCCrHCoV2pfBxwIkqOYw3oxt9Mvl89+Rsv
A1Q8QPoVMHNEDwKhdZXzPeRdmA/WB1/kB0lEwXAjsUz53bvV+b9x0nILQ/FKoHaS
lAjlDwuLwPxdIQc7DX7ffAx8abcTJ9RC/z+POEvgWlUyEHC54k9vobghN41i++Ur
8cbRHPLQ4DR2kCB4oVt/IIPgq2pQ+YqQrBXRGw8/fYR/ug+bKBdMY3tTXbEqpGXk
OL8PgsE7tNOdvDO3jwVdHkNS/7OZRCdY4vyvMtWsDvTCleQvNbu7+fp+PaOF8Ey5
LOlVn3t/NvD4DaeXNhI4tv8brSQP6fKHjxCmWajNCl/qb3ZcEOBNqtLpe/hix2fZ
3ca4HrG4yXW7C9fZLskUDSF4rFEi9xn3gLbkv9rqvOjD7KNZG1j4p/F9hxG4EjqF
Uf2Lxf8jMJBXUkczPlIiGcDGCqWqN5onzHUIUVz/AN1wlQTNIAQfyWxUIGPXv+cY
FwdroNWlYqskGtDGPhsCoGBg7oUDSjd7yFj+WPEL1lFTuLKN0o3zX5bBY9fMHm9h
hyqJHjIugKSZnkU0Sf0CuDOobLQFD8l3aQ6c7y2GOwDPv5N8McK9Y5uCY9IW6XXb
U2lqkQzt+xKRH4xn3SqxTBrnxr5chej6Y2pP/d6SkwurHOXb9h4WNHHqMWQxsnJ6
HEztJdwRsm81t35cKrbGuR75KdbsRBlKBOTspHI2miguCik2UyOXH46CUKUS1KQx
K5SAZqMikhq0Ppou4XDwMcuVOTtnpHDJ84VGqN36kwN+sTN2rT697rv0VDB6Vc5i
J1lpBiAFsQQVPgb1Nfkk07jjuPXTuEEVWySogmiO2bHK20qadRcKwy9ufs9kSfOS
EYh2f7hOOfHAGhgabJgY5d7EV2eq+keLyueLg3LVifmfqbf4uTs67ZPX21YpmdOV
4m3Rqh57LQkswngd+jnMrN6yWXLUl+SGEqd/G2nMQLeoUHAGHDqRJB27IdfK++0M
/Cp8cIi/FJ8MWDS2BthKDqPyx4GGrRt9n0uB3t5WUDOBE79+RxuAN2pzOMBMXKal
0lkOuX2Pfc6iw9r56COuwmMSvd5yHOzGpRNKZhP4HCJt5AJhjI6HdFIWjsx4d0SD
7onC2kCPw+KErx2oJxQ7q0RkP5RR+CrhBb2whagx48B7H2CfhLSBfPDaVHIM/Xox
vmsU6gI6CbtoqNnMVz2KxVGO5ZQZyPh6ie1lndEHsvxDfPbX1Vwr5lsPYyPcHQ8U
Qf4DMKzkk+rtM85q0YJ+1K8JHlNafVoB/RBrCHeuaupkqcSQrXNdcDdx6ablvRbU
eH6kpRsYzDOAUcjCXjfTYQs7YcG+sBRyAmkzOPWwW8jpK18uoEvaGmbjlgrU8zui
JpU6YmY07/c61QAlUyC/j7JjwhIfMQ8LNNTc/s0r7oSq2J5adttDa+XGDBPUbSnE
wuHEHXdmwvZVsmbcH9ZDlPzs8Qf/BNSzCYn24cae2/ujHChn+qGXqQXKMKYSv4+A
jQr7i5qalAqYcxB4ke6ROolW/YtZBMq9K3lSYs9LgswMT/Es2r8UI4lkpWoqCvOS
eN4WPJhzpl1AQTItQJ/a9R9RUxN+1emPr2gxaIfHNxVQdLXHgRKQbVFJdm6hYogF
Wmvq2//RpjtzIWBiWpRvFayGyTHm0KE1EugJjHBKIQUg0In2OFzQWy6skdtQ7LA2
haTbpCEVXsIVRP4UhvS428cPi2V9idBIthXIZOVVp1bpStiJgfXNthT7nsXzXCcq
vKjqpIHa35oM+XCIVyqgBg2wFq5C4WGz5Qr3DX0ysYoej2jrEUdnwlk1LNJnOvnC
dzZ+Np2hMrjIGyf5+0EUB3ECIclYTIc085BKWIgTVnwVxZCcjF37cn0zalmyqbjp
tMfsaQENDX4LXHNqJ1SZG58otMuaax9k8ZCiz6kr8q3yYpaFBIyGGASZG/YrrO8A
TcC0dDl5g6Jo4jLqbEGh7GZgpgX3efKnx7LrgTX9Gu4WEWm7ns1cUSgVm5AQPP6J
srK+FMhLhDDjZWdUoWz4JZtVQc5pRnoNKUKTLoT4+RPK7ke763qhTHpXC4KSTD3k
va9cOUDAnBxf4MTQqXUvKHuDDO232S7y3gF8WD3rA+QAZ3FV3FCNnLnNB8s7dwRa
8sPn5rWCD+oqnE0b35Y3zlZ3TWX11wtBgqAUS8dVQaxHOz5M2JIYM7VKY/e8EJhW
eShwzhhnmrBxQCvXSNIEH44hAgaLiuATiqI0BGbIov4DB9Qzet1PnJPG7jHgpWYo
oe5mhRmdlKDIcekQR1K9co2dwGfwgYR2urjXPZWQOfxNAEA4goaDKqfGMY0/TUqc
+n20A81bZJ2q1JVEEne4gIr5IGAhD8rzYELx3K/ZtZKn0nG75rs/v4bfg3YRXhri
ER24iBzfudCPWS0Lb+EAzE32GUWUj3A09pNxmSGbT3l7AVcQPdXHRfTwQckYXHkb
96LVYFPDmCgKsSFUGBQW7u4cdt6u08cdtGS3/Ch0qvKIriwsNzILydxsBE8jJkE0
NKCe4NaLv+GWWFfutlm3Q7TY5gcB32YcpJYslC1jsrk4+hznoYhmYHoN18V5wdbY
7Ogw01fg1HCc1LPGRlnY6PwZGy/1qB7FOg58X81BkFMOrAgmyLiN+N7Q5gvYZ7wv
G2SOQldH8qzOnjABpgCtkZtbGx6GzGB5jyWxjIDDrjUAXov5oSTNKynymjkb1dVK
LMFDteqeEJVwvU/iebwH7A==
`protect END_PROTECTED
