`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48kty23gjzPX6QVlml+UHGbxGP/Y4+e8UVy7eAj4uaTl
BMlL/+mLGhGADQ14PPv/2f2SxMbw1iKUPJxi0t5Cqxvl7ed1wiEady35OCBcgbfT
9jnlxzrsEoBea95zPtfZxHHswdObv8bO76hIrvYfS8P0uBV2be6MG5Vz32pCLIV9
lMAEAcXNZzNFfiHhpSl58UT1G/yRbLNs/gsVZ1lZ5DshvBabIyZ5OwC1Cw7q3OHE
DtQJVxrvzcvn25aPH+2NV/UgMpxtmZ9tQFneR3bMvWykgZBoG8cS0n/arG9Xs3/m
G8w6J8QBwTYxQwZLCA8ZGw==
`protect END_PROTECTED
