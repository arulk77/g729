`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
G1sGRCv4XY0+ZYKAmhCuAtt6vAdldEY0Y48U7qEFv2T3mYco9yLQxtI1unj6kTJe
J8Pna8rnZgcv5vFn8gj/Cacw7hqFF22oI1dyUP9QITFq2FRV7q83pgnpGZXMFY5r
YxYN3sThfLhFxD3Gxf5pvIprkkJrZprhOBbbuoOOrlg=
`protect END_PROTECTED
