`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SYdX/dZH7vUxU4QVaFij2lg6uXqel37rxdZ0F0z9dpe4
2lSdxhRiZEaicf8EPFLVY+bIlyIWB195wmTc6z9d0B6yjpWuORX2qX/emArmdf6e
3wHNxpM6cb48DXH/k9MgSWMwsX5BPWgslWSepBloZXhJrgW7ogpzZRS8o46mqzBd
2EkR2OTixLmJZ1a536jNVmveN7/bKU6+xBt4Rhr04WTHeARFJRWV4Nb3d26UBymu
ZuA9yHC/5VZKCbGlWuLuUdbpv9sHtrkbZGlejgtm8OubppxZzEvs4E++648Je0ov
K1G9jnw4P2xJremHQN3b7f7RLEubQmjvObIh1PtFBZJA0ZOI2YjF/4st1XH+qWXl
7xZyy+XP5z1iXKguJTIkP7Wj/Led79fAjrgsxeHaIyciKAvk8u0FrvGrTuQDghJV
nCCIuytMP3YRwQnmFxIpaX1FeO/f0VCD9mObAqECiRcn/YQp415VcxcDWukxsw10
b1L4vlfoePlb8NQ9TnofamDcW0RduZPpc/MbbjKnAydxeoucn/Og+XEBy3+O5uRG
XyWd3A8LwCRfT2reCveo+7AfGvqZc9GSyg3hRhy3dn/vOmTwBUZfU8ZOdiPM2hGO
sK4WKnRKbbwOaRShlZeYmUahvy3jU1Yh45rCu33Nz/4tGSJnzdwzx6YoRMXyKxJE
sfzf6xP5sPPoj/yrzDfP1AzI0TyUZSAP59s1UkikHH7NBtjAr9gyOwnDUqUMxm7o
aXdTUHjXQkGolZd1q62CrFbR/mB2/x/0IBT8h1EjferWzDaOHYDp7noLAHaANZem
`protect END_PROTECTED
