`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QsjRDfPuOD3UHvxlNqV2rquL/uvu6NDKSOk+rgOTwNNFOMs8hQzoTF99D1onmnmj
kyXpUVY5Yp6ML7U1B6xOqxGL0AsXmJYwEFHvOEeGD2wQBNzY5/Zut25UgXl0+E+L
vgvCxzQ3eGqaO4iaOejC5syVbTxNTKG7Dv8ZZGir4q1FuuScsp7FnAz2c4A1bWX3
botTS0UELPaULGONC2LR3mKw6Cu03QEG5W9drOsLgStQXoE0E90Jyv6KdWUe0tEm
2qzMRoBXi6Ygs9gdfRD8ZKHIV2/cizfl8wkM4xFGttk=
`protect END_PROTECTED
