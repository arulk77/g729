`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKl6hCflltVZZB+H4gn0vWhM7JSQWGU/iHMWwbMjDx7d
SCCpyWw9Rd+Qhl2HTHxMA3NoF78lV8LY9ZuEMlME03sEqDmrk3/eCY2ukaXDV6fO
DXVD3H8iMJrND+dhYK2JmZK1Bud+xlJXJ9nYBJJAOIj5DqzmE7DIElYZqC+1ThAa
Rr4UBwSIgzA1rmhjbuIuHlIhUCF4+2f9co/VCSgwbEur39ofZRjg6A/cK5zo53I0
ty1/jQlsjKCXGqN3ayjlun2GdBvJg0izu3QzcmiEztL7hyTrHdKNkwCjD8xDzXkN
E203GQw0sseWs6DzISLwAcR8XkfJwF/RtGe75mHt2oxDGOuNVzi9xIyiLHVwV64n
8L7QIdx3e0I76n0fV4EC/Q==
`protect END_PROTECTED
