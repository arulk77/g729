`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAd23gNT5zo+30vp5jLC98aDI4X23FiXLVybTB62QVSUP
WTH7qmBSfVoZ5PDmS2ok92cpJzkz4BLmXKh6P1ZM0U46sljcyzGWMyEfFj29s5uD
GywDk+2ADAeWjmhbKxXBqkBFojlSDxkxeEoBh4lgm+TREbL+91+hOhseGtKakzE5
Q/mg2U9SMGyXBxLsV8/+CC/mcWbebsUrIclNewI50DMgFYb69V2xIRLCaVZocWFt
Gpi7BQStuqOY6LmdPRmlFMGXrWWDzFpvguLRuVbaD/GlI9LB7juwtYTk8fDOXJDJ
Lbif18rTquJusZB8X6BNcM02kvEt7+F1k5hH55xZLq5kyhvP5pfVZJkPx+rn90Hx
tDlfCNSu6Z+cqHGM0HHTv1w7A9bdo2g0PyZSK5T8Wr5jpAsO5CR/4U1uAr66Ieku
xGhCSUcw+1dw56j6Cp1pfRa77Ke5hmc5UT646J5PcsVaHSziKsxeeitX1CWPtQlW
2GbSbE7hvtqvHrk0j6iWnYvsYfxWixNWvBg0llxebS3VTAgZJmovF6z0qp5ndfB+
Eb8BgyMU94dYNnEn/GTepBBIvpcRdW/TQpAlQW5eDJqjtCG9NXnHeRhCULlpJYpE
aa/pVU66mTvF57EIQL/B3nn6qQ+pOJzJyeQLQBcNDu2Ef4MP3HZlaXda+QjfDVPc
TFU4Zjb/M+ogrhHj3K4CjOc4b/LNIwB45x95oYoDs6DpY8RK+SaUfEi3jgzy8CID
bFV0kg2fLmWJDRinz3RiJqzFEhIqIisvxL2R+KuV4iflevHIKeGLbztmBGfXF7Vf
Ia+h0rmOKNyuMep70O2zyUDiaR3qNI3DVnaKPTQFzSL3Ff+vw6bBMTsE/pYUWUSN
UyFivDkf3akcHrFpi+bKes6RSl/VOJxjxWWVxSsNfXcUlpA1cviljR2RI1UtZLI+
5oXjYy5VZMFO2HoZNCkFzf0q4D3b5vbTg+1oKV+WHg3ujeIiQwOt+oqHP8u4qHPZ
pOXjV9G3MaVU73rDiRU/3rEGawxZpTGCroNPH1+2I8qaCP0gulJtr9ga3DsL1dDY
hOVst3q24IX/9euDuaUugXzBBO7Su6qbIxnmQzScYFaK1WiqT4sGbIcGfQp170Kj
tviHHLY/Q4fynYlEbCY8jlWbUqoGFmMLD5WNUfhptQWg4dX2LASsIG2axHLG0es9
RV1Idf9ELyAGKbe6SBuRcMmUq0FaZcgd/yRrJu5L1Lg33QbTU2Po08XNMfXF+6cv
aYLmNETpTU5ORqOCAjF/0XV6J7jGJBEn+NmdkjL8S05ElsGoyoUDoY6/5PItsizT
2eAkkB0YkR8rXQHN7QRCabVyEXGE9omKx3WyZvCzhvODwtXa8d1OWrWO+l7LjAea
b7F1W1OVntlU93+CKNprZbnxFpw7Dt4qmoBuWKGg59HmvT+7xyGP2NnZts0pEOEK
+JKDsbtvNReO9tl8z97Asw6JYruh6zakyLFbeAf4VagR5FGI56yt+aPslWZ+rMl0
NgHlEGba5mGftM2hoa5rSpZfohO+GX8ErRPDFar+ESCb43omRquc1TJfOm+YVVlS
Bc0HGxlSaWBRTFcjH6QmmCV10voboVXFzKgqocsMctpI4tyazO9eo8U0lJHoOokk
pGmFnDaMuHChj2R8gXewof3XBHuNarnMTlZBRBR7wVNYslDGTA9dufctFwS4JS62
82T3tTJJ4RsvCJ6csLxyTBUhVl6Pz9WzUl5qNRqXRzhcgS/KVmaUM5hlDlq1/1/x
6bFm4aDnUOra6jtv8YFwqN8uWIfSG/ndnNY914IuWtImIJcuVUrJlMzDKMlTsf4m
7FrjrM8Q4z1a/TnVQfxXkPWvsTmneTw1nSNjQMSxVBA1Vy2THl+I/uAmDFJPExTI
a82tt02wRuQCSK3Az53gP+subBK8P9H4TBfVx2cn356GgjIZ4tbyANnSIzMkqPrE
qgn+G3Yce1ar5+jKypLjeKwsQwWO8X1BvRtRpKBS8RwrvHz3AbPQsNCJ4TnFwdCd
XiU55j9PH0nwYdCUubCJXiEqbcYmhXYyeh7ubKIYkYv4H5aa/3DkZXXJ1WZWgBFu
qzGBJaUqrjfkQFQn+shyU0iLy7UnsADKumpBXK7lRXlQv1fuZ5sr2yNJf53iO35j
WcGw6YkVLXEmVEQ8bLm0Az7/WEcsLG+LtUdApbTQbIlvs1+rY24K32n5zZ/yPwc8
YBcnMdxM3LYfusuaixmFtFYNSjVKoInIZ9Xd575Vvj3Ag3PtAreW/66/iK9+o/Hk
dvAVecdMRCEprB8/d8YyGQnKecsN/Y7lpGHDfN17X7szfrSVm+E+GLfq/Bp/icdC
wMp7X1jaMi2qPsqYJx3gIliXV7M2fUsjUC3JUH1pitjlNvjPT9k9NTmpdZz33eG7
mRWSeL1o/TSMlewIfQyt5cl48DkxsCQmkM6Ptq13L9sElo+Q4elzXncc0wutKCQ9
2On+bYfU00wHpg8yxHPYOMeeKgHf9KbfHibXKejAsleEzCJh/x7pWtG8cce4Kw2i
Y5SHfSQom/l/T95Ip3LOr1Ill/nF47aIr1/bOFWq8+BrUW5jUA4a/OAwEWVggy9Z
g3zOm+1IRKWziUbWwc13Y/gBQ2LhsbeG6qRudYNDbGTIcPe7SeObrvZjlkjSFHHb
4VnygRqw418gFz9sbm66uGiPbUKWcYff9jLtZRLaEY6z7mEGaweig4lOEtFh7yTW
lIAsuuJrwEqemyAVix1z6B/0yM6sPwY7cv3L50Hlpj7M5Tfiv7u4lLm2sTh5uD10
npI951l1QxWr5oQI/S4HIMoNlg/D4fTQJPsYdDazCCisinVeOujBkrxLjtYMQtdH
FVXV9ZQJ34VzWvlWUcVTPJlYMQgvKI0JzOm42B8+0EIPhG5ieRAX//rRYpmN0+Fy
Ptupj0GSd+VsDGBJ9Q+lU0CkGvEpC9NBuc5WelETR0RtHJwxQEKw6YMu4PtJLVmL
kYKcNdiHfjRlDjBHAk10f38xnRg5reBTgDdLmZrXxmkY99o3eC1qifCP0wHEZXN8
e5B7ydb9IIYHqTz1PQO+7mieTYMX8UofcUnAIGsmn7ydFM5QwDnwwJwhk6KQQPoG
uRe9dLgrWembp3/Lc7Eclw+cBvUFSZYUxhx7BQi4KjDWiOrjlnlKrI1GHNoUxPde
FRGXPs930WDOxhazKHuwirpttYK1trlszSmZ2RTdAEnSoaXtOMFO2mrJdqpVGMg0
i6PnDsfiUPoSmdDq6QInM12VHxjkGOYoJv70WqJSZbwu9QYTTl9qGxRvD9o2bb6b
2bDtLx2mA64bBxTjJCYIJPl0A5+Sw/9Tqxt5bFElkCr4BlPTsALVa9FhudxpkoMp
f7bMwLtlduyWwnFwhJwyncUPeR0xn994HIYhXeTb5XUK2giExZ+BQkpjtvQ9FxDh
MiKRgOr9ANiv3zEl9OWJFnyp30cJWxjUf2r45OVybEw2NwDAhXgz93QwpUwD3BX8
q2nP0Tb4iQ1YmgUUClP9XKoZNzLJC4VkRYJvdWPwY4ei0JmhqRfKgfhk/dcrXGdH
rv2LlLVF/umUBsOKM3s6ZenyP35kiFrED/UYNQ5BNImZnKKxUIltVyNG+x9sLtFe
RXoys55gHxCX6Vc0D81RNghpGMdilNSOgC6LrXK13JhVzSWS1jNrN6LpuVkkmO8M
HVqVg+g5gXglZ7K/S+PFvlLBaF3dNWUUJkbgWQs7nR/ort/sCCR/WnodJe0wDg0m
k+VlTHEtEHgxio1yjr2CyAkZb/UFXsdsB9oFAxcAcYTTyuEFmvF6+SdDRY3XCKJn
OlXCEzqdt6XfR3xY1SVeC9QfMkLW3xlg7Xr7PRvttb4X+1xuUwv1rIDiJtOJvMT/
3LAj/vpR0VuWpy2Sljh8lYASKi0b18+aBT4wGZA0/Nl0sVJIBN/V1R7kH6u7yxk5
SuWztMa86+UISR8XxVLkqirM3rnLPXJtlSBCAWwAf4SUvHxYjnYh7muHTvelZCZo
ZSqTOfCtsG1oM4ITlxKktV2MJ86HrwADssKQ2Q1upqONlzrisTNj6yfNaLdbdi0F
qoeiiCZIkUzEqN9HUI7jvAoQ6ITkPmnvB6rYNOVEM7JZtkdgTy4cBayDMdvFk56S
5zawpsXQBYK8cJOrGx/INT2nS/7/bUNDpjDeBcDR0qey3EM/QOZLT5LRWVeB8Xr/
IClgE2hqw4JAobHo7ZMyEIu3UuY+4sSVYN0a7qbs3X8lglwwV+m5DAWBRmCSqOtF
jNGCpCZsb8xBstJoALCIxmDi3J7rOyYjr0pePFID9pn+rqA8MqR4cmWkyuOXe5Nq
X+5SpCJlrS5+HpxQkOiQvVTxiilY1Uw+Qe3hGqUkVeM1hM8/1WWN930VXWfbiqWH
4xNnLhYfLXR98LPW5Tasl9BQMG02FYd+YC+Ds+WkDdURbbOgX+xV9Rq0LgaFCINU
3WTnfo78WtPvx6jYiq5lEc4Q3o3w/KJTu1zneMUar4xFI5sPmLKoL4tCfCBTog7t
nd/C7AsPF3nM/Rm/f2JIKmZXA7GnHdr5eRx9aROvpK3uRnqJ8fL452+izaey11cM
JZ0i/e7xzlcZXftXgJD7QpPXsLRhljbyhYv8qQtA6uUVnVOvGgS3nndkIPm7pVWM
VW3d4/DgDfUiNd3V62ixgQpv9VOpD2R4pNzUgD4dNYX+gPCN1QS6JhgytcjnnhAK
Jvz1fDX9DZJ6A118sRRUf+sJU1YcYf3hUyFMFkdImkCceh6W4RumqCEKJTZ25D4v
ZR51m/Qr3iyvKnmqh63Ti+hb5WGFVo9dlSEAN2LbIqAIx5QyQMOhF5gz3ifn6stF
eVfmzkowIbydwJYp/72Cs5fTprc5EqI8iTe0EBOzeezgc68cqPqCOeR4lIi5EZLg
B/HNtD2Oi/++raKcvBW5Q2xaIRtz2gTuCth5+4uRdrg0s6bfI2UX87fRM8vOM310
4nvq/711AVlfcbMzuAqLIonHQ7QR4md0w7t7cN8eWon8jq84k2UhDzF2EsYhbz5T
9uQO6J1rVmYrtNlfdE0SR1KM58D4V/SN9VpwiO4Uys+1/H4s0LmFKFbAsl2avQA1
Vw53Mvkul6hgZDSxBAhs2iMdK5W5mKwEvUhg0AOH1jevbEuNgqgbaa6gh4UDwCa3
5t0XTwAHaFlDDeSKR5RrH+4gxgNO88eE6ijGTAd31CnAS5G14/M3gO0R8v6KBXSG
K7ZllYIbJlXGXoMYdvEZewdYLjZeGIwD1SkDdO4ys3zCdQS6g5AuvPgOitisbT/4
qJNnNOVmfG/HHTWAXQMiXkH69D8aRjGItTbdrR6fh3wZ8jmUhRE36ohpkcoh//hs
pQgRbtI9/j6uY8uevVDSbUDU/BQMr0rfvjbDY3EVUM5Sqp7Y2zcaT4mDl0YX8Agm
ANYKAUC5jkL8c9PqXx1hncD2uYGV44/48Z07vwiy1FnEwoMNVhfebHMPBw8qv0jk
eZzHMG5UJ3/lNatcRBNF0TRwwaT2CnUORVjSo75mv1ljKQ/MuqxVWMOm4MFEG5WO
RWlPXDhdgzij9tmZoUIpEJ4ygG7nfkj33/92HdxqAWX4tc39cPb/YTV08Q/ZGL4x
tZdV7UYYs6os7bmzdxAICZQwHi96HI/qgtvk80KsXdskRvbRvqYk4cfr63EDYlMS
Xct525IqttNeA1LVCKVjsE1wobIO8vjaK4hM9uJos1UVIquCZpx+djMkz0NpiHF/
wVKa7/0hYPYeaIIgwo2HOYpef+HivG/dL/aOK3944HHYLHlEN2jk+06vqpT4O/SX
wSMrUc+VVtVTbmfk4K0o6GtqOk2R4YpQ/5e1EdJkEaMey6guJSvnTt604WFyCmWs
N9SatAa9hf9QFlug28JHT+hyyAR29dtx4L9tR59v1lAIAlMAVSrm17T1EOuq3hjf
9xA7wAlfpVZ11InI5hJJc+m34GbT+OVOWPa0/Mh6u+EwsT0P1hZ/2Z332leEh9GG
zfcHmQpkWv0tDq10qfwlHQbhZJA7V7GXWyOmnVVcGYJc09eLuc3RywuffefRNsPU
q64vMf7d20CK/+Q4LpXylGXVSTcRojfXV5KwGah1J1tFnG/Cvk0WbTo5YsiAgwiL
7BRFcXSx+utihOofUMnfVsYrKRBEe8bjOQo7R6fc7ovuWcZuxFVtSsBvEwT0OTyn
7k+Dr5oEYSlWhuStmdYr7wgFDTKpqxFd/yiEqof7ALPLt7wxfH/KUXlztflQmWxK
KfkFoWaslkekrzUJupR5D1xn67lAO2BUE1UQ1jR+Q7re7QFlTgivNVStDAYaVY06
ynsKU7I+S1CohUKQuA4TizIVdE7lGpneuagOlhIrgXjAeZpLH2LIf0jyGnyZZtY6
7VARQNv//h3vOeBfpzgu6cca+9zeTCvtEu+ClJFyUxppcewn8p3Mbtvz6ryOKQxV
23g9gWJeTZzQg2B6SKACLieVlyrlBz150no+9rQCkQ2kqgdB/ESCcUXtuJxpouTM
I96NRAWDfcjd2ON+FvJ0MhTDu02+1X2rJZDhtVDbQH9bHCfhdKZLoQa/uW7+Xyp2
ppZqCPpn4c2Ktk/UnJEuCpR4shFBAK2GBtw8qoHm2RYSOhQtBmj5sI16cjuShp+B
lRsiveK7BAwtYZ2IawTk4mIUXol4X0Pb9dZr0JvcP23osxDj8YF53V+1K+pqbRqC
0J3rhk6cueRL/tX6R17F1VQN7wpp1iumS38v8XEFKrb4vqD2LEgwtb1OKWQubQ0l
jQ9wnXWanIchOoyTDS25yJfomUq34yeFxNme0S25z9DN4YwbGUyMOcOpnq4UBbKG
bskax3EF/3mKsLgVeH1FOTQf/pTXnZ/fzd+UtcbnTc0xVCz90ceiWVVR2pTsJ4g/
gg1NMS5cu/9o3xa8IB+gZQYAg1gntASiAmrNGbMmIAF77uyGEmB5ILPCHhwfPjfN
2l9t9wLG/Ek6WzRZnkHrnoRF42D3Y5L/LeuCmPgflJ7e6+mkOdEpnx6hBnSienNw
NMUcz5GNfmyNoP75qD8vhMG+F8QZ+Y5JuZTXbGYU1Tsyz6tyewoEfEStYRBwF+VY
H7/keFqg2bwwJUa35Evq0MjGApogGyDItTCA2lL5xDVBQV1CZ2wOnXufwXfoQcDp
Dw0/8SVIUMESeec5FU7JcQtLJcXGa8xRzKh9McoYbINheu00GTY9XwKq0LiXW4aO
zREPfapR9Nxw77wt2SnqZixvWEr0rzI6S9fJGcQA4bO/U7wVaRPJjC1aqa0mlJaA
IsCC1FJM3xPOO+WC+PafVJTPtBmgNrn2B2xWFLPeIlVpL562DaxKNuopFgZp5AOM
4hOfKY0paQ6TmCRZCaNgBexeFUDmd5+4+Yh4JHYnVbr06zUWjso72H9B/VOlvDr8
raPXh7GubkyT3XRw4F/x7wvtAnlyhBL3o1Li93jA9L+vYkHnYEzTBRPVlOfN5brN
tlsIlNAtQyL36FnVk7+sGLD0LNwba8sM9YCAA0eYjjSbFqLtqcVZdtVh4pFf8bWy
APl4thf///c2jkk+fyPQpiCpqsC9w5xhYN+yvi4r2h6DGbClllk3LGEG5SQRgvTQ
rT3cg2RoGRInQ6CyDsf1x06e0izX0wnP17Nt9r5Mz6Pf5xCfAO2gKzKumTsmh5Kg
qIIssT1CK2dNZjwyjAU2B9JInff038F7/1W9iGTb9FUq+n7YM5m78a4B0hEirssD
pGo/0wveWDePM+N73eagX2BYp8+MAZ2S/0qOmW1skzS/0mXvoznpKcvw5BGU+AKO
p2VxUGNZMG5WdV3WQNTIgSvMmMpBnsTBl7Ce8Jt/XZsVwwuThWcm1iZmXlvd6v1J
pSC0OWgwcst52G52wqJzN5YTgyWjAa8sus0WTuxG6FsqTLUKWo+OGPBfo+IedaH2
veU8oxAn5fYyQ4wSQ7zrY8DLchNO+VakULvWGyMtm1N9WHi+MRUu+E0w5Q1V7eWC
l6LPvfGv/K55bfuOBVJUZEEEPOL9VC2bxnt2V93W3uo5xC08H//mqkRubAP/69j7
DbdqKyIkXdk9njAkD8asKkLcZSUiK1EIm1f7Gr8eAKEIIVTPwp2E1DpXVrJ7lDYa
ZKf1SFr+LoESZC67uB3CK5+hCNCvAJRS1+URAAPQooP5X46ll/Ma/NPFc0SkZyIx
IJHaHF6+Yj+bweqaMKWNDWwSfFNrCcvF8RJ8Lj4HqsBCZTywcvS/lOMXghSBWMjd
G0wYSzsucXhzLUdPYrTZ0WXfocb6MgYcdlZr8PYl4Dfx9G0CwYuAl1jBdkvDC5gL
om9v+o01KhVAVxZiXXvRq6Yo92vlo6XywAvzp5d5UxPb5MUHCYbs2dcSvzsmfJde
ZPFVbTpMrXnoq64wiNsFoj88v+91Gh6NA6IGZHBSep2A42f9STUpzf3Tddnmk7/5
jzB0CJ0lOxTyJ+an/F7tciARqQMtvhL32HwKhySB7THxiw6EA5R/2Ld8Xo/SX4Eh
kDz8pkUOhxRL74X8yIeDR4A9iX8HaEQqF5b/2a8D7V9NTA11H6cxuia43Gy5y/9p
PvKcPTMT2BQt9kmiL91OEMhZajonIKC5UonU0IMMvD98b99uWGJ68oEfV4BEARCp
WBVs16Zf2M1qvy25xazhzeUZXToGJSBjWxqr9gpnoK2N3Vur0NchORf1fKTM0Wqc
Yybf4t0Xn1PgG0vSyYgntgCqvuKXy6nUh5yhUgTDTIDVkthFw63wuh2ZKE66T3cD
xB4cvIHq0R9Uj0+h2GFxdxANok6shkVzWkS4iSFiu73qeDYRKNZQN3rc94hwixVz
S7NdN8ENTO4fC6nU/A1InhszB/SkXTdi6ckSH09bdOTy/gvF7YjgF1MEM3Kmzg8d
vKCELgZ5SJAAykh9pvCFoWGwVpG+ZqzimqDNtZXtry5Y0nb8VA/BllJ4whHU1102
Ch+UQ5plxdB0lL7eJ8DEp3sigckcU3rZYcUdrtDSS58gDDvsxugWq12PSJIcwl+d
JoSodb8elNxa45Bjae8fZf/PYa8x6dmz/GJ0Y9HY83eX6UV6giY58jJLawX9E7RE
oObMqsGlPflJxR4XBqiLeX4MAUbt9tWUFKKxskf4QYPGjXHVsblyXOOKiQila404
Jb8xK2xKRIjgsDTFpxO5bEbeIzIvgVEHMjnrJXVQgtivgSytrU+uNUx6T6W3tlUc
XTcEwvtyKpXs7pVwE5bu/ndNWOfNjhawKirnTMwS/gY2daSDNzYjElKbCPDc3bf3
be5IIjmEBzSHBtPZJL9kSRtnC3hGYS4WulApr3eoh0w2vVEUfA4DZIPGAiJLqglo
rQeWkSrZD1K8sKBAdv1G7KRhbVHizc4njnSWFD0ZFY+7IVWLleotFondf+9WGxxx
yefdJlGhbpZzvZKwVghq+d+qr5694Jsy6KSUwQXyCEOqvxHqDUV7Dm4Z/g2urlfx
E+HeDmiqF3dFSvAeIXf6xM057c+bHw7zMlVf3uQfs0bUXYpqQwkF6UKa1WIKreFn
+IHSWl7RT8515E1y8Pcwc+AiRwqNJck4bJ3o6FKKch4VSY+xHpQiIFHBjeMhs2HW
GRRD9hQrFPlnmsvkG6RsKVQedk12Vp0vcEvAVYOq8wSlD6037PsOiAyhp+DaTa53
FJe5HQuaBBHwYjDKHXdD9y7k021Nz1pQ7nig0YFfuRSPe8/31PjgbMLIu7MuHBPE
dct4054sW9OFv6gc4wMtcqnwUKp8UtJgWf/DjylggSUlr4isMUB9VFi24OT3JFgX
lsSSLp6l0PHZJJsr2jUAIIrAvxu3c3XOLAD3S9bHXz5/Qh1qdmyxlhT9t9MKfwX2
A3ds8JQTmYorCuccxC4KHdGdpq05hApZNmLqThy+PqxcnEZ6E/rPFn/GEnCze1G1
CX0sgDAyrw6XndOFgL0xf5yFWvNNY6uviTafq+usymeDVv518fLaQ+hpWu7SffMv
+ysT8hMg/BFmssU2sYeISDXFjJQYG5NkTP0JJNBBhrTrtmlNp1NIwTAkZhKYwPK0
7xJg+L0HJrX/HOkLC2Tetij725hzgHq+KTaVXkEiXLWepl33ZDpKV0I4W/sAVaG6
53h93qY0NtYKlbzTdx7cmLII8CEUKZAyRaAcjmW5pV2Ophax2DD4yM1+YXLKRiVG
b3hUKkpN5pmPWg4+IF4m/J0gdu39FmgXjOJpZAzSCbusTxDZMW9ibCleyr2kAb5a
Qm3qHPR3sZ21AzFsekTZCGn9Hilt8XAyK83KFJEHtKGujpEnjfmZqL+JZYre7JEI
IMm0nlkCaUUm5yuXNfCBDjCp4WP+VQPItqTdgJ5B59cS4JEc/XQk2+phWoAZ02+U
yeuDawPP2yk3avEs1H+n9M+6tgFK6zuMSCWhYoTqsDWoShrmg2cryQnCfhqzJ6UB
JjjdR3BsP7lvLcgxoEzF8T6VnYwLjWpeikWdF1WILel4YahqdumTdZ8DXZzRtB2n
LyEtgxU0HwhKnnx8F51Rx8IUtDWXnWYSCbZD8MLzYHcYPXYroSdXMjuPv2lEiCup
zAvQvDVvN7b0tvbuFq9u08+O/o/oFxePv2h6I7rAp6QnoFJrGcUOFOST4YfrouL/
QmhNHd1sXsZjTFPEHnDBqWH4JNaO5QPxqLhVBQWEcu1ZENOiJxr1Y75wRn1kXUW/
nUNBIRJhN1yf+hH0aEdxA7+3qdImwAdU65dMewQiSG+BWl44F/xRCRwyczxPvsdI
dDHupyhORssYFe6bIUmgCH17IFAy4DFv/NmkPgGbagnBIsS/U3xxTLL2g7jxSw5T
WK63pB1xYrD8YGYtD+w7ppQztPC5/G8css5+HQKl9rS70GI/8qGDzUL3+GGzu8sR
kjRfd2M2XV1KU2LBJ0ekdsyAXn8NVHuF98f4Yugx2RuyiWziYHuAFurdGiW0r1cJ
Iwo7kE0Oqzuojnywzv2U8xGMGPJfvyI+m6wyzbmj6WzqM2rqLcuVWmr4oyHzIqmb
k8sn0Ixf4wYgenvDRYxeGHcdJ1i7/LwPL0wPsEd0sQ7DHIx5goiKNC4sE7vpM089
18AVkIr62yZtWHNWUmEbbg6/shqAQQjncqISaZ/E3U43qswN4B2VdXeom3KKkArj
YB98q1Jr7gNhY3iPCuAYeXBEZc3uD6/xBN5xo6Aa94+A8EvoH5cQbB3k9O7nSsQJ
x5eAhQrP3M+5B3JOGUxZxbWis7zMMyyv424w4yRS14PBegbA7+nLC1hhxdHQ5xKh
aNOgaL3rhO4LiDt5etgqVLkccVE+2BH12doi2GBPw8m6pVUqKd/BiP/GgTwZXBS1
4wz/IubXkTcEQBHpswyDoLbLtJpa984G4VsAVnlhtrerBo1Mn5T3s8zQxxj0Rb28
7CXnCPi2RUWnZTIpNGMYfZ0qpo/W33fN5g8gqtl9gmnydxZUgan658E61ZIeRvNM
+4UoybeX86QowsE0fLtsXASVdhh7h+nEBQ2huupTPvCr3hBIH0VAGZmQtBPHkfxF
zpz315tTIM1SjV3+LrNdEfGKXdFQPj1li+W2nWPv1EJNrnlC/CGMRKhgprzQSAX+
dqa1fyVWXIWqMI4k/f4zpzYVScpRXv32XtBKvmqxMN0xnND3wbIakO5jORWydb88
TZoYtTKr4vnvZCF4W6JIvwIC83FPEuvfyQC4I1+knoWUKoxfz3LH95YaJhhOVU6/
yE9BARmCWniiL2VuCH5/01oGnKtehUH2/Q2bAd8G2F58Dd+6H/oFfZvDtU9VWNPM
+u9ec5zPfeyUvclXlA+uV5mc8j7DVvFY/cigS5vs9XOm+lNmeTkl375LMw4vOH+/
IE2ezW09qtYg/n+vCY3VCm37D8WZv5KeqIgcfUr5fFZbOHHfMpUm8fUFw0spW5Ih
xMel9+etyVM/kSkfOKSh4v8zfOnHfU197fyUJksvEZPiGB1Ok3Fwivm8z6OAGKb1
QfxJN61dLTu8ANVZx0NCfrtKRWI1wiTShfEr3z29NhWf/Wtp3nqcEXNe3NjEBBMM
a1hZARoZQXe1I4QSqbEiZQc6v1coS4lPY1XExmsl/hZqzDdffa6m4GKOuF4CkXwH
u1m2uI3R3v5BVazvDYH5k/SKWbs+9X0uouY5sdSwHRc7pa1p7dy/lg1HvlyDzYkK
Hrhr5vRKerVLmoAuScMnZtUvQ5WG2d84dGpO/Hf7xSWSL4BeQVPQlnVQW0tiLvJK
Gm+/jn7ve9xsPS2/nhbk60J8cRqfGXIPHE+44TsLzypK4YLyy/uUol0ZZmFJygFx
CYOfsUAw82PZgf8uRZVYZNvxqQgUtoBe7FjfjLT+04tO7Z5mr20dDcH3ijhaon+P
c+suKhVZzeXPhrXaMctKIY6V4ACGLlbmSW/6/800ricthePt1NgzN0SIwVKIlDfL
3DdkM6VdOIf6vt7MKqPjQdDvJs8VctXN8Shu6fDL5/fEJHlxDJrmdjB/ZPKeJ1oD
xcHZWFayO01oCVjLVjfahimCJeyzNh++3MMYnusWq0X5DjHu+i1xhiemeFc4veQm
2VuqE+6efJsxSZhSrf9dBH2xt28ShpoCJAGYAHeets/clIRZULsCvj4lGow/1ts4
W2J+MEYv0v9esaMshq8Ci9W9HM7BloE9LwcV2YyHAUcj1+f83MqVj5MR34f48Pd+
gl1JTCHWsO5hkGi9GOVoMm+O5HnUOJ8J6pG0zNBaLu/xKby0sO7PofZWXqg/QpAP
4zee2aXraQLLwceSdl89MC3u0+RY+AbT5epw8KSRhoEF9lAEvL4PMviXmuNV28gS
BWXdl0e9/GztP9n2TUfkVizJ2g68nuql/b9xWO0Yav+2LcKKqJWS9HtWIjhkJAih
rxNqcEKiP5LmMlwsimpve1UOZU4mr1vSSCpVcnISIZXMiwSlv4fTIj11J4e+3MPP
4bfpOpT15Hmoo/Hj8fRMKGdTDd4gE3miKKkR+9wWTHKRueG+WAcELBOw4vey9TvU
q9goqXQntlQaCKNawOFLN5hvamGFmzdD5hAiuftL1yej0drEmR0JE8qtOwmPHDlH
qQ6/gKTima8mO5pKFMVshE2qDJfvKXxkUDB5fd9kW2aXIY0VbBs4Q6rQiNiwXu2T
yNl6ZtOktsDo5gOkAZU7ADWKXUM/g9h86aTksKxMCaMbt3E4Wp4qv3Sun5Ir/ez8
zPA7fNMxHj8RWddeMXHHd8l3TwVT0cZpexv1PbhgsRfHEik0xsRU+96+QNjrBS/Y
azognq2gDmYGao9LrTqFD6rpuYGgXAI7NTxtuAt72gdEZrz52zGXHQtX0su+TGGy
h8QEL95P4N45H2lVw0ex9sOY7IFN18KXQ/f48WsuF2WUfejlDOwnQH5PPZeYNc8B
wtqzx/A+5Hiv9CvAu+pHxyZc/M3X5ksqcgL1ge22em/N04yyLOB4064omW5NKIgU
zahSVi0VQspJj0EXDvg6J3G5Eh72dKK0h8KVri15bFFoyQA4DZiUwBbPWeS1wuhj
al1w2lXnM/VNmL5dwKXz9ZCoc/inTWazUo8TVSJdutc5IJBbWgYDVLogdvNHK+DF
lkk+NwCe2gkjIfjnIFI+WvCp2RjpdrPXKesRilYJZMkuhsoKCqQFtFnNkPbNhGHT
rXiU5WmRSDKuINu1BpeS8PCgZhI4IG6y1srZ1QjdHZ0GZoX/VSwJAIVx8f74gE/N
CPjWgRlow7VHQ0LQB9QNKf0URaljWiYK+pvvfGxZLNo=
`protect END_PROTECTED
