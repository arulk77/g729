`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGMWH6AaQYcIoxGcbdMEHC4LHgq9FbXjIRNPob27lgP3
/8hWpXeycpIwb1k4FciVt7XrWTKdOnGKqIFeUavcVZihnN6+ap63bSNIzklHaJNE
R49pmZF255IkoZaiTE5nAEUzuvQFJbEaG3hP3vemP2QhtwpKYMTpY9bHUBOKFyxz
X+7mTuVh/mQClzMG79GNy2gEsTDcWSQWwyPbw/qH/YQqAyXppN24g2TEkMrH7lS3
ov0k1AGB3QOZJNoaOzUBtN2JW4HNqzTOWDaYf+TtvfK9AWDaPJmraRyoWyD4XUYg
`protect END_PROTECTED
