`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCA0p6yuScbF22gG/cL6dFSPpBTfzrmyM+tpIwJ8dne0
OYwqHHdhPoWuW1x71wQ+oBSH/lzdAd4GHIDxWdOfiLzaxMU55CIhoN42I9u+cgKU
2F6m6BlNwxuyNW2YwnjfCYwMoZIh8SwE2C3V7gRraEUxfu6RXP5sT1LvlG7H7bgG
oFUnY5mInDbEPEHBQ9Vhtm1LIAiG1OlYM/lQzvY1jFqbxoD8pXiNA52UcIGwnbeM
vETxatG0NQRbdExOtaru1KanRe2qrqQNfKMZZ7VMvuzs8gRUEs4JqxRx7LTZN0ao
`protect END_PROTECTED
