`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DTuxsHB0qyMswer+vvP9FBmmstFG7LZbCelladxNQ58P4v+JVYtrUbtTN8Z/KxqS
lx1z6I925+rP/aVX+8jZRfiRmIkfgDuCS3TP1xmomSBFSOtmwakGyCKpr43D1KvW
C64lmaHZDwFtVI7jzAB9v4qzU7mJguUJjJeYAoOscb5/T4W2cEAqUzv7svu1RikQ
feoANWWpBeZf6kBQqFCfrsXQlDWUiGR38QBDXKCQed2/ZoEespxB7Y6JzR0lwMto
dR7Pgaa/dsKLVU3uB79N9blCK+b6O0FohktH/l7VoJcreItLRjBXHyZ2Qfnn3C/O
aAwkq2PDcIpndc+dqwauIfXZUYtzaoSzkxUJhotiD8c=
`protect END_PROTECTED
