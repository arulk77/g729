`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOZn4rgjk4VTQ05s7In5dPdApsolcub8Ijci/jM5OI/f
jok5kVpX6aBNnJ42lBQslMRbGcpR7+FhfLnK0reBVePj6y69KeCGUUrqdzqHRRUv
Bw0cz0gdpmq62aIhrixYG6VDf3me4o5eKyiXLGea/ivEf58CrVJ/jbitTG8BKuAB
XFB/CGgmBIWlcLrJeWmXB4OpeCzh2XcCykcAJOkle5U8rL0wa4d6aX64kjUTXoyZ
uPCj0wZAxA/qjrTUn6oQEyzNqu4ONTyZTwbXh2gV11ZVSeTS5w4jhcMvxpDcMHht
bH3N3w4fN5yCRFJMNQ1wKQ==
`protect END_PROTECTED
