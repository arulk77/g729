`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C2Kqqob7nSHAGW5U9wiTc7OAPtWPp8nNQ0hOv8qePo5N
dBxoq7qb9DUxciJbtBrnOdViypWy2hz2CtzHRz61szJdMRXQo3I3mLX6dlTDDv4g
4NULzRsQjYKPblX2AhaeJDhHYvaKF0/QJvF9P8oFnNrWHpHKohGBTdOIRH9ioS7f
xSe3vRUKUjczLx5UYr7qdNf9kiLH2GOo3P09qHdMwQV58JO92IpxymW7WDvGI7VO
txLtju+40i4zsM4L0/ZvRs/H67Uaprbgn7zzadq1StGUMqXKVdov3guPZLnF/vpv
fpcQWEIUOTfjNa3KrDfzrqPy6bB5WwgZpALw3Xf1wbM+F/l6BlYrIB/FWY5JPZux
nyNauQwKtbnSB6LUypOhF87CVWZ5QJHVA+Y3xAX52LWvtvovtNlD+D1qKGKIP76N
sXR07V0OcJ9FmBwMj6t6pFJFf9JiM7m5otExo77I0JxofIMJ3ta6Z/XII2dHz58u
DFpulzhN/1JV1+Mtz/ni814x9B92ExuuS5scwP02dy1+abf/n6Q2sXCotvYg+ic7
`protect END_PROTECTED
