`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA5+oVmdvjiSCbb9sabtmKD0Vzg2HDC2n4VllI2FyHGJ
VloOYSeLpxHfuphUN5je4tNCoZJcPWDbZJrAJNrOczIj4j2lrTp06Sfvm+1fOwzv
y7iW141wtpImjMWfF9lV1AJpalu3B4h3dxEhhhbg4XR4kBrXckSt7NpGfj+J0e9b
Vgp12pKY9CBZMgiRso62UBppm/HKjswu5+4X6kaUpSw6MjQInCifa5YyO1SB1rlB
grrRqHTISyUswuiEizvZr4vd2pNJiOkIOLIvL7cI/JOQKsEL051/lXa5MVJpXJqF
/qA5HVJKLnjvZvhviJdkYJdUImqaKx1mfIYHknH67iTni+myq4cFWxZ7FUAuq7Ds
`protect END_PROTECTED
