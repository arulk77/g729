`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+g+4qEkGP1mtrYYImSy6xWBG8xkjYxedReFfVbBE8gk
8GAljGzvOAJTZAhnYpk4lWJcNPvpehlUwE7ItggHauq0SQrkRe3up+iYgJNoTpqY
UrtYTbcvfSAptuYaW133TQv0LHuNADi1fzFIB2ou1lut8OnQqf9G1B9d2TqkpOYn
P1yclSnj83AyeNEXSihLk76GH3DnIS/K5ETihDIQSRc=
`protect END_PROTECTED
