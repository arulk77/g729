`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zjMAXuZwZikPFVi9vqHw3X9C32RW5euQCxEwQyVBtHn
0LlCx6JeyVXKfhotTHdsVfckRPggIiZOYAElQE7TqitZYVy4RF3ZP6Yyjhw4MgAk
IonggI55VKtSuhCmW5fYUrMJZxuFrmjXjJiqo9aLQ8pQQtYwiqwma0i9xiTviiXv
kOqaIX/bI8aT5M22Wi82uGCFXSbmmzNB61jcvgrigSk=
`protect END_PROTECTED
