`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8TxMo8bFwoRinC9We4ZhIB15Mb8rJGAfteU2J7kW8qQ
0Cowg8RTIOH2bk91DV0jexv8cITciipMl7kbR22mM84IlCjZeQ3fX/at0lji/9sm
939Hn7Ve9apoQe3dU4AjEinWkaavuyv4DijuoYAdMkilL3iT1K1PTbPjBYdh4oAX
IXiUucrMT8uYWWKUnZqkJV9mohT+TpawGWRPgQVd8SuQUVR28dzTdddgHKKVaa0S
HzI+lPiHd5bKWCGDG42nJlH0dlWrsSrBGxZtPPGrhOvXehsSi4NFHsCmA8AUJqTG
W10zVcHGlJyrYRVBILNr/meJncOoJ91MjJM4Euq3xLTFprH5kBHuXciX3WdXE/BG
TIGCEYiEv9x7ZMeTGtIFGjsVpqeTZJdTUoion7Y/5acGzVT/qSwo+q8QAlnEmqhX
SpzahR/kaPKpcbyhhMYf6TA0Th4qH7S69L2bnQXYwJyb2KegYWLLgri1+gGV4dSC
TM0S+baUnyNh9L5uoylggH0QQU/gxGS6Oek7yM3c/vvaMk+lJfN/gdwwMJFdmyex
QdYqzJ14gGUj4CPA8WP4heE4y7IhlDZQU65FYbbIt73ApZPx7T5l36Sc6xp2wUQP
HchzQuGnu8MQ8HC0ThmGYk1eArOG3o0qr3z7Y1lp8rLRc4trjHPRSNRLGpvjhmjG
ta6XB5XQgW/Dth3oJeiKC5nj5mB9CA4ICpU8otNQ5YZ3lwbYYga13fGgkQp78iqm
5cWGVm7FgNZze9xPVYQfrjh9oXnMB+H7dRsJoRwHtL7PvG4374zEry5q3ZMnO5T8
VHt0WEReldYrKi+02xQkt9tkNqqSmcakPEB6Xx1TyHo+UO4HSNQrm0mPJZUyCsjr
p3x/3yoVzUAurBja3nDxep9IXfcdc/UxlYiv4XYC/XBikMjp8o1KCQl0EGw5Dvty
hBKqaI77ZXYheH3wdFq7OIhIDBeg+3TS3BZlqpcMWcsyTbneptMpzIOPCnrod+JH
3+nuq0q15NCSR9m9MtJ7rd5kHPL3jzbF2BQBb+pByKhElBj09z8Y7/86b3MzIHHJ
1G47TvdR9OTd+Or8pkQShEuc7jv77ix5IvB9BFieizT72QbEh487AZf1MDUrgEQ1
nGRsFSvkP2VkSWZ7KzgNPb54sfPrX4YwEYQKlECXnVFMivLPJubwLXgNya7xCcDL
wnLBZCZt2gTIAGExpW9bG3Z0JLBPO/fL1hbMfWEqm7gWvfMxBhO/nGxUtdpV/lw+
B67IL2Z0G/x5fT2xf5eAQue5FKJARSmeaTZNg4j9LknmWWzyT3D/9U1HMJEVQ8lP
6nR2Iap1PynVTrf8zBOs6xCeyNyrK9EyHM8/PJ03Wtv6OhzpunH0sWfmcLLHaddd
OTn+C8J5tOBER2/Bx04wkW+KCBPwGsbadogsBMAmV/lEPM0qbs5F9lfwRzCyPN3W
7o9fOtC1g16oH0ObNyRBC7kr31yU6bD2fjP91ZffFw+BOUVsprTOMuFxDpp+mK21
xwNzCM+2+QITqqyaTny5db/gRYNbwnNuaHAespHhix6huBTSlJFi0KzcKEYjsdGn
+fzxyBw7ylqOXLgsG1jHcPiRFkbU7GWalNGEyLDTBYXvyxLbYBgQi1q628c7YVBr
+q6+GNHQobS3r0uQoI5GQsFe6e5vDYK5GjesYG+I7Ndr9s8QjqL4Ee9iSCEprnWP
+HqFjUwm7OVXVNpCy7sPKoGEzp6Aih7awgM51mjRWQB8/gvPJjAyGsIOioIYEzhu
1ioMUDi5OkbIs6XAo4BmSgwI2PsK45WTlLpBbF6r0UoHqpwAKavT23cOceBgcpKc
juL6PrawLjtAYmUakunmbodinsC6GosJR0njZVphLyJEV8uY9UzqkVvhgj6V6y3R
CEi6IdYVifl8wHbl8wy7YgQEUN+qwH1hT3Tqm5YeeoVGJbfSa8FirXR9tJaw8o+g
7f/07TaG48P/5xGbx9zhBK4Hj0jstXwX46Q+hREoQi53gQsCzMULiShZgm/1F8Mj
9iFCcwBQvrU1hAXLPDoypG2S0O4CkVR8Qu+2f2cbOBzE9m/7sR5WISLNB/878G+t
i9bFsmhlap/sIWbW2YIRwOKSDJLLgmX6117C1jMXXoPAPMq3iuUFsj/1gFkxq4xv
uwL9sEqq/7qY0aiuvaGA1voTZ/Lq+nzd7LziI5SahhnBsrR28LUo7vefW07aL4oS
3UHY8LxdTBUivyNlYhictMqyN7CgFfbvTt3iux7yG7TYXcTd+dA7OMCqbDrv/hl4
aTQmBZb+rW2mnua5KSGLVLx3BGdWVS7Dhj9EM76g06nXzb9btzPymg4LORGc9yo3
0R7BQaKD4YDIjILZORENm7QvnaDPRZ4mvlJSZ7qZi0VrGmhbxgjgxR0e16Gv/Eb1
mB1C1ygVZS3M1xM3Vm1uyml1J3K0yHz6SmC9X4uNuIetM1KJM6k9GZs4X8h53zWA
OBmL68eOg+cbMvv5OwHfH2CX7+2Ln2unHOP/qOsb3fLfLZHAWZ8JBq5sEy80BPFq
RpqjuG5sJJhz8lIy4opG7dXM4Dsm742s8aQp7chYWm1zTk9DPlVWlvB85IswwVyQ
C+KmSHAdaZ4uus2zZ/Ygt/mMFXWRrMEWC43ByTUMcCHCXi2GFdbdnzFcLkWQKlqr
f0fSgVEkaRzb6rhgsePkGo+RiMjG6wS9hr+RucFGnfZOHpJc4xfxmZdgE45kyh8G
qdJEA40O7buDblXWbvGR/ZThStAaNOaYHe5EkgRabKWeTfDQt/AEVTXjt8QEvZYW
70OS1zxRbKWdaUWdastVuTwmR8aSTxeDgONTXuXTQMS+re47IlTBow/RdxoRm2DJ
Ncj6JLk1+f4Omq5YLEfwI/8ZL0+cLjizc2lZDtsifgzGsol99c8uaMybcx8pq2n8
CMD01CoKs0KE4uvKXslDh4HnogU+zi1FLzK3qbsH62beFDH8R5HcjCynSXcKOsMV
i7XYzzJ8WlBpnnWJVHtD+VZEXhg82swllWOdG9qztePO7PSFj5Uo8or/3OlOy+wy
SU0B6FfCVg2inAOSauh9iur3zbNtmVzSM7+zetiWwlbz60LmCm5kbGzrWMMQQypj
5mP9SQ6sUpruy+eil2oMFjvW3rkzgUkDNmMlaKnFbkxTR9xtRzoqSaQeyqq/Fd4C
20sOr8GxGtjXs9l7JVQDDrFasSuLzU1jCYTDUyWSO1s4pzrt2PHTNwO/fPnAEcUQ
8EUdEDhBH/z92v2qIqmEVbY1JQmyjisbxdLuuuRyh0Ef1iKLZWJQ2SImRvkzPSYP
2NMGBieMhrB1qH2LX/nNfVO8hMCxWJfguaGGeffaJI3EKutEh5TNjpKvCwPc6GlB
pdP4sWuKLSAf6Bm2hVLdOF9np0t+uXX5CCej+QosmTYeM3UN6SGsIOQrTrlU8XFa
vPNr8s3UOD9KwWuBfiN5eJx1ucXrR8wWvq9bBCdrBkQ3/4U5jk31xYdPGVweqrDN
0PI4BaZVa2+01w9ou/4mtBNlEttkwDWEUKy7mJ9wzstggf5xNafV4olW5fcZXeah
JZdmk+7EX/6FQ7Z/TENxOsq5LQgCMTHFiMaJRmJnLADJT9/NeH+3tm2zzDD4eoWJ
n5+0aeaxnyhWdYegwLZZ9RMzhlRtEy/qCPva1/+3OQOWzOOwgFC1yMqfZvjBpaXE
hCce1QapBnkihMMn4KxnBkd5ZqjsdUvUoCHbk7QUubIMKt2DVtWo7PQ05bsia+LQ
1QfbvTjSPOfJe0/6cxxTRrBTRo2lUe3QyouPcP9rJYtSfYioMojrZJdSVFwt5Yor
awcgvtg7H/FUWuBueSdt1Qztt/BhSywfFgJVm1CkJw3OOSw+dVTC/aNx0B6C+Mqa
HMBwvpuX4+bcGHlLTlStOv4XnfhknqvAeMeFWYTUOfr2SybdQojcXauM1Gf8Fxzv
TMRajKEIAqQsxDCQnztzPPp+T3320Jyt4gUrN0d3XwQyPBvF5XObfYwyoLNcdbs4
XgLDVSVqXFRxqwOFz0xp+ZTADx4cvZFSD/I5g5Rc/o0JfmicljjjFKkSuEE/KKqY
XLH9M7KGa9Ymy/dom8nurNMrzfaIbIHpw3IFyBTZZue0Wl47UYg5whlrXPZRcNBN
KqCekZQ0/uY26GZl4MVQWbOeeZiOmvfefhmyYh/duYJdH4VLxXIL6iutGK8zAGrh
RcYGk+sKcE58bhRQzWNfwpn+ei9UTEcyDDXPh9lGF1F+x5YwjqIGultYWy0wq/KS
4rWMrB8GdDgluOrVqVjgAbrvoU6DXIzJarIWc+dy08frk7OQYbCAdw/Eh1V2rq5k
wAUb9Zd9UoGfMxDePtiUeko/QCiU37dZeqASzZrHml9gAwJcEnHe+rvD5WUNYOJB
BO+wpUEZRMjgPLTZC5xAfVcOcB0tGw6qhxZXzckxmkmv2L4YgXmU7uqL2jWx/sDX
PHAP36RbK+PQyaJu+8NBN2yTKrCUwfMO2K8qMX9APKEUEG2mtamus4R2fDbsdbVm
KQtb/n2F+r2PlzwhQMs3lEfffN3CadLyfyel3UUXc7PiuOPBZe8c/bittcDl8wbT
45GvebzlScoRk29/7TXNeBhN9rTAHRGGRK2wJcFyr1IpTta/W2E3VTFNpmwpNCxp
2tVQv6i8/ypNIDwNrknMTipyrXtcyk+QG/Qk9HTiXukhhgxC8bXj8mETJdMeyzjI
DdshxHOvi2SKDUA+CJ/HwCvNYU8b1CwsE1cdpm4KLAB50s5Lvt5uxNzWAKOyH6Ve
dLCPfNUZsrnKwFh+BG2fHJD8LwbEHJy/VXV0o3EKeFnO6HggMcH5n4fm0F82eFRd
naJfhlg8KAXEbiFMz9Dn3196yXi1b5A73TsjC+E5Ia+oaZKfJisCdLtB7zLA5SZP
VQeaI1XcRZ/AKt/xWA/6A6/8WTC88AzXrn4UbrMvsIYr2JWuTRDp9RaUV5KZA/1j
HKDpsC5njr17jt8IySxKlGn3bKpKwcreqUYoaZYL9iM4MwHallFOWmfcw8iBdusR
r1ZpV/H55c5/mZFjM09vhpkjB/YlVRpw5YG0ENMVIqH7xr0STOSWM/MVEva3YMPc
gKbU3idFnv+8fD+XBIhbunAp1E44hYQUNXi+yOV43DOncy9VpacjbTAzeH6skKow
Rafwdu3iQUjdIFAfQ5f27Azw07lMSk25p/omatqjWCmUvpJ+XxdmSUP1yEpMTCu6
Lmpw56pT2qyRsMWwrHTn+q0E5DHPi0zvN5yH7pwzamZIRG2UPAYtmjiTxcoeVjBi
mlBQIplEk42AzwV4dDBqgQYXvUu6Ms78fMZ91jsqwYzhA0DliYFkUHAcaKpWnJL5
KFA+Ca6126bhgWNyGb9d+rudBJoJwPGJY/6jwFDdPbTIO4aiYnEmQ1aPtQB/1YU+
UQjt7u3wptQwJTJlW3PeTC8p8fnVQuiizjyN8MPWdS2vb2I41lp2dxnHFjXtbl1c
vc8xgYWQJehxdcdSeLppeoiQaanQjQc7C3UfX4PbosaIUbgWaG57DP0ETPtbUug1
/fnO5CNifTPo8/uVwGH+AwpXV7zKMG+5jJfHYxrTWpRbYxQoV1qufg6SBTBV1yoY
CXlLE9i/KvrZ4PhxMMD3Au7jH7XoHS3SmMavmb+blzccmNH82GOYRvgFV7Mu1SuL
JMSHX8DV9uXWgXzG4/kwRUj6t1tFtZzQ/7IxSABRFEthaz+LGOM+r6qsUYse4rzb
HCnvVcKfPr2EqtpEkIbiyIrRIbgvGh0LBfKnn0eKJxoLym51xH7UFJZo2zFThZii
TH/UbB/QYIGJDxDF27kAkgTVp2/xj5KVwBEeOEQAO15BT5HgPASCb+JUMcL4Eaea
cTZPaly4LFjMZwwx1c2RInG1qUYVa95lYJaJ+5WC5BiZcGG96GNIhOkUMa4OwbRQ
PLm63hsIiuoJZLMt1fRRBX+bFFh4wEkHY07IMNGa0TSwQFSIfLD2kzXRwZUP5WzI
72okEzjQhpYD1JLhK0YJ7zkky/yWyPt1s44TCdx+0KhzOHF6h8i0Aqy3Kva9VHkI
JXwZhQEG1rWCQODOqb4XEIj3AoUP95zsx+ekeVIsL85OWREzrICen3FI739+Dbze
rzzj75lTz+L/Txlps9cc5joM2qSNEenBraHUhL0EeebMri7WJLfbShaPwTAOo+mH
l43MT2ci57TR53wmnlOgx0wo/7DkvE8eVNI6qPCPMOdZbfNxuEfbmKhv64pooAB5
tDTMjAftD+5xltMj684PRdyi5wKvrJdmm1ZZjnZJ3DjNRZEPS50lTcMstZM3aIlt
q8rURUWbQ1yw/PLj2zw5fySDZGLu0sdvABxnuc2rARkNrwnQumAp92k9+fGZ+Qcz
0fvxa0RNgeG/FJ+ymDUDgxkD9U7f62npRcGRPqzoLyReyp0z29dkqTKvVQhYqA87
rWBZdla6GFGXIeCbWjZu+JBAzmP9iquGtPdTAjUt6rh657vO/h4XHBHnRN2RUigb
ycJ2rGTb5M6M6jE0KSafnXb/IlqrI6uxU4TM0dpdZy5RJzoS1GzYpZJse+uL++jc
fS6sSLA65iW8pLMXUlE6b1DjWAsV2rJHohz0mtftG2SIB/jD8AqpwSR4JRPzG/lo
6Fqgn3KuGzCmoRf+v+M2EijV6xKlQeoBGx2zkbofyT2ui1FpKrVU4SGm7qNBkvBp
cGSQiDgyKtkkQsf3koi7zofw0EL952sKD9sghunIe+jus2Tgov2soysUrx+VsDip
wFtzhe8PIOMHXLVZAMNtEDCnHC29H/1jGnEypdoyxHvSUg0hg2oI7u1UzAA2mCO1
hV/oMg7Kn3DZRxzSezKbxqRCC1QWchh93zmqRJ8cmpc5iSUhFHIci8+/bKGx2hWj
htoj4yWZB/+clSVLNHakTAVzMmoPa6TOWaca1YHHFnxM3zBW5ddo13298G8GIRRs
1nRfKfoq98O+lWDnTUrzcrt+baqqLg3SCcigJtcbVfTUgrEW3Hz9mmb68UFXYjJc
l36aLnVvxdj2pCfHQpQF5KuViKGuE7APBrW9gzkzZ3i5zmE4cTrRdmTiVXekSmpf
9D6+NiwUyQDFiZ/mWrlDzgoPQb+PX7Dq9b0hKjsP4ivthBx3wLm/t3ljfAT2u5Q/
9ituQNs0qBVv1ivBsCWQJlrPg12WgiKuicSM4AXTwWgP50fMB/VDmcYtFFzpcEs1
NGNKmSv5bddnaqb651QK7LvlYwLBSiwVk8RwuHSkb5yvTQNS4s98fK1O3hEK/bY5
yw83qaSy7vlwiGhfmmKBwnkEdIjgxuTImQcBalpzUmtyLClPGG0csK5fFCHpHyZu
+YyvknrIp3/0lU5RdFo7PMajnMfwqivlH/NKiWwRBUL+LqCP/Gav77wFk0WWGBfN
SOiJwaq5saNbmVYBRWFuBytTmXhQy/2GT0JmA9z/xLymAJsGsZt3WrGaCfxMd3kG
J8mbir8KTN6ZEPM+CYF2VQNkAzeBlz00t/9J65VbfH5qPkRJIYrI8G6NAyQ9FRpz
XZS+H4b2GmKMcr0kokuAZ4b0VgVFIXMoCEcb7fq68zRvGDuWSrOESnmx60O6nGij
O8mY4rSbuizYzoU3ySG58SvIiCW3VVIxnZ/LOIxyflEJyzl6FQ+VmboUdGsFkzYO
eVT3i8DwNuP34SoV0wsUdZ9Dbi9hwKfTW6ln2CDAz7e98e5HXFqI3wjqVHLG5whK
rtR7TeKj47THtGIfKA0KUjHHURWkVx620VWpr/UM11r3t1LHaHzrMqO0lpEneZa6
CTU9mtlO1FApvCb6+GuDG+uozSgsmWpq8J0hSI/j3K67xrr99Y/5AoafnC3zwY4C
B4eacrsYj0X84i6QA36MZXa0Ed0LpLHlIp5ZdOawjng6IKBlg/73v4AAeTV4cEfZ
WGGqowUlCcVC86e4jBqnNnqXpNHGrys65bg1LMS7+X3hpnjXa3UIgTBSubyQwyBb
4wb1M0dOxpNBlmv83csqSZLoJRAN54kb79OGNrEdvTdc5wTOCCDl0aJcUseDtp/a
AC6LOLJ5upa1fXTQf3NnbqT1cIriLrLmmZ4seIOHCZFrNbV1EvbwQhK8CQ3dqdUI
n9sPuDhV5iiBRJD1mWqT0QGR7893orMJKooyTBUzkCiSfKe3wO37FAAbKkIOolxv
P6yLMYbiL/P1i0t7/7JL6CFpOru3a4fHgjvvWkHcRTDu/U9hMheiGC2WFrPZr6VJ
zhWNAfBIjilpW7bwoW5iZ3+oPka7otL5T/C5Cqu9mAhy0peIkcqreU/FpykKWvt6
ul0nSjc67ptCyjWlFSc0IeSPqghyRaLeO12+SF/RXq12gyrrdSaMTch82Uav/1ki
GoifXHAA5on8hYhgKvlLbFoN3fj//JC7J78zRcWlZlqGv9ruQexnGj53EzDB8CxW
f4MR+/fSYrg/n6cb9e+XSi+nW9T2NULCYat5/qI1VQDun9RO2vy5tWZZsGZUVf77
TzNFZ/QY2zjAigqMtitdf3UU/Swk45XKqLyw5I43hOd9f91FIrjay8dgBhGPeKxO
cfpAHG+af94SN8mg7/+4dbOc348jQ5SHZea9LEMdPmF/fUily7Fr1fGedUsNS/eB
+DQEp9KrHfyf1DkdZ4Vj+4u7szn9LvjsR/gp9tCy36BTtC4pMLCIp71SP3Pg3HA0
dDd1J/MQUINeND44RPmIP8QGIjEz3BAWXBb1O4EPzRWhrT4+l+u4uiN9A2nM6yH/
aCuVKAXZ4VkbJVWpVGA+k5zsmMU/GoaIIlfmCQvl+VS/gAqY9GzDGGmM/hm1FAxR
l2YsZDFuKsjq00ydrd+lRJP66GZjR5YLRs66I1s+UN0SwXxwmx3TNYT3YzVVSC+S
384CicUHoarsG9unjDXN7rz+jQ84URYnXp/bqkVfYAk=
`protect END_PROTECTED
