`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yCC88EXmpvwSeRGLgmPWuWOw2GY/KnxOwTIP3hHVRyl
wycqk/8bVgNzFJ59ANHVX/ZCKl26PHwLuDvB8+PHSbArt/fNQnMnhbm9mkcsxvp1
rD0Xh2l+BgokLcrpzdLqrips94+Z+3d8YpNPS0dC/jEpHiitpoJdz3UWfiQuoQTt
NNl21+vIbdGqWi7Y4zlWchCjYwHCvT2GoNfsnCaT0bygUWG9W60FLqmtSQZloQ/0
Nx1jKDp59r3L0ARaMfoJH4KIUX7tsd8B8Eb41blXszzcGqoyFlbcjjSbD8j7sxN8
sbgvNUnaLRvSj1u9WWt5bswD2C9E8QvTJI08tvwfjANPv9Z/Zi29CuXEhmgRk3fI
HLQocQdsBVkY6Tp9rcOXRA==
`protect END_PROTECTED
