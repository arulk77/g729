`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFZM6w2OchIVYLK17DqrcpNYHk7Yion9GhZ9dd5xxNcB
Cz5Q/nqhA1vDUUCtm2zwuykqdnyDW6pxqqnc9KfHGm+i7RXBR3ez1fWBVbbE1Uzq
BEjLEO3M26dazE7hUQQJLxOMoBHRnJOekjncoEKIiSSpPSx2b//x0otUNhGaL5LV
yj6BJCPPOzaeqlpdpiDu+83ILzm+5ymMl7pF/9iP/IuA4WpRnen4eWYz2ZMd4BLQ
zlUHueh3m748kxxbJ3jd9Npgs7quMIGxJJVnF/A+NzO2X5/Q1CTEnB2Lql7BRv7I
dHQ2uFOtcuLvNJpnepNW4NahBsyOO809l+Hru2GGi1UTvfoaLlfFBsoh2EvQRRcc
rK325o5qjkEsnDe8DLgYUklN6EK9AMOyJHxdobfVfF9Yj4z9T9sMADhO5RAhtRW9
rQ62LL91HPL4nzsaoezpY2RwO4b9k8d2P5noBbuOCUR6WejMOW23qCndZoluNWTa
kxF7QB0sNF7n3HNGF1fR6Ez7M3NmYuIMBdTTnYWfg/LdsATglV6MU9S9NhihqJMd
kyV5zk1fBwrNjZyN0H7at0n6aRyVa/aRj6QXn7h3pGsyCsqBoHg3b7fe6n8AUFzo
`protect END_PROTECTED
