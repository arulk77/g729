`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAFsuF85fpM9xmydrf0WRQiY5QPwrr/JN+dXOc8zFkAy
cT5lrq69/P5AG2A3d7PX/vinohScCNF9maHVssK32DSWZra5Y1raDcXiLMy45pZg
dN8nQ1CATkJUXNzjiorlknNwXLrK0cuN7mW6BBpZpDV3lsbPzS/NlhMb3Q2IUTDl
9ZLY+UopXA8KkfS0KU0TN35DQdiT7kPEpwNhowbWhcW6o8812AkXzQcJ6ZLiSW6W
`protect END_PROTECTED
