`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH9SrK90Bh8iscdZLY8B0Q58e1J+3j5NJupZ37MOio1w
Grpg6W4z1OCTbs3eZKVc/f0RI9TxBN4V7aM9dtePJwKW60gqlF6dFSDqme8ezIk3
DB3xL9A8rLv5jZi3/AcA1C1IvfTKjgOW/aO4jTU0BJjb2DD7qVFaPVPWVcxA+1FM
jytqnbbNXoNuALg7Sn9N3zWcQMz6Jes4S8eiL85BnbIwmDi8Wdyek5GIzgY2R/o6
DQPXeUe9sBqdYc8O326mwfuEGe/x2uR01rKEyKOWkS62REJSrnCwxTsssRnYEQNo
zRbBTOjMTjG9SHnA16BHk8LCAulhHbog/YQHBSKon233Kgg9KB6Twb+Ay4IahBpk
DP+/MMk7BocL35lkiktIe3PitTqyX7QeWdyv8cMsiy8f7RmcAr3OumGJdvHmUGjn
BaUkZpw619cZok/9Fbbn4qgiKhWGsUNtIwABkJfgc42icDc4C7jg+LO1tO169XWJ
03c020I8PB1nizx3cUYBepu2Kc1dj765Dm95fboa06wMIIO7Z6x13C11kVd7tRue
KwGYOeiAI/mGh/kpglvtkqPiXYiQW0jtEZmOFSyGRE0zmCpXFp1KbsPyvVvr2+yJ
JEkv3RaTNQwWfvpY69MePkW6iy4H+4jDepamihaI813QKI+BYtUgeheaYTMM21jz
`protect END_PROTECTED
