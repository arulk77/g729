`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAPQzvVG3V+9ogjpWGPbrIJftDIbzPo9+hRChqNqTc1j
Gd8xc8VNv+NkEX9OBy7y1FuodTXVUVBhRZwYLhDF8sDINFbfP5yY1pI+CpyEMGVm
cc243ejPS3T3EdEvKFtBmnPBbkrrAfX0DLehBxEUYyI1+81X8r556sUJbRXNULDa
s7PuETrnsocs6ELhQ2CfVynNaUToRuhlkN80e78lE0bn0yX5+Qr6BrvVEgHi9N6F
X0TlS1rG/mnCpkesyJu4OySho+TZLAeUTH0G1lPKgOgPzYUTbmeyqIut1O9bzOyD
tjvdnMeRXAoUAiiGdPjfZyWOjsp183rE+93BUQ8+U9m+S17Vz5qHuukH8n9B7Ue/
XZJi4mf6xHGXwLwUIjiiyKCNAo0ZGM5HQRfzPbLFnP11cNFZzAcpfjCf1qUiFblK
zJIVbBoC702lrGELFZ7UOid3/dUa+ueKjKmZW70u4JE=
`protect END_PROTECTED
