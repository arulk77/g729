`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aYbyzd5U5aA2oJxe98CKWydDCUTSMgFpqP9WBt++b80e
Aeqq2pgIzmzBSf4HlXTmrl9s5t45TpD01ZOr88jpjsU88KpwKs4Fq8Nxmmaqr3zy
4ZhZku9QozZNbqjv6yEZApcQ32aKzOe4cnQLHFawrLYK+3gTF16Kyvlt6GaI4Hf1
8xkcxbTRrfy58dIxKUewBldkBZ1Ls8LNWGbCSv7XMa6i7jaTu5ySjQx9b3RewO4q
/IxubKg1jLF39T4dR0wDnJRBD3/iY4ojeQFrUk9A4xMsugG0qMx3oUoz6VJB2RRL
`protect END_PROTECTED
