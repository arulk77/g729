`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C+Hb5Gta4kh8zOkRNMNS3K32DJNoApmlMOfTsF0erjvQ
dW34EuyY+Hqpl0dR40DipLvwDhAc1FhbmPU4bycBpjoVsoEGpQYxaKVuTZxJBevu
yxfEMmHk77avw7mIAUtMmctWL1+ZFeBB8e049b7c57wClaaED+k+HsVe2JP8HAWi
F8TCG+bKQZX9/k2YyGfn+kY5BVoczz6mLdxH1Fk+zgBR5wmsy75Khwasok/TwFso
zvrxSW9Xt9E9ShbvZ+oJPG89VcwyXpJ9qNLrtj7w0038SdW87RrGmFU9295Y4f31
sE9JoU7+3/9SKTIYDaV1NXhDl8fHg648SWyD/po8QLKE0T6rl9FtaeZdFfnclYxq
s/zxZTbvtEqvCLvwrHYADUy+S1HSXVqoS5fgG/eXzZ2nHU2SKyQeWu0TRRoF/E0C
Vg0ku7KEosBfc8VEFH9kFvPFPsIxW0UUNxWECx+yOCS46IvjDUrJeIiS5QT4z/iO
E1p0XcjIyLoqAqzoHr+TLIHEoiUKw5jl9iCsbMVbd1rgZRvbCK8X4scNwTT9M117
9OTfJzWmMef7xb2hYyTjKKD0/trL0RNZIbE7J8aAS8E0NCduUwF2dmHuHzUjULNV
eFCtoD8iYATZlFVjOZphO2r/KOwbl5WKmCWIA7vZ1JjuO+mZpCnD8sa42BtgBAxO
kJv2GbQYvLUdfvz5BXswIIUrR9VR9/d+NydFXEDqoPm8zFHhu+9mBSM8KPdjLMzw
5EswXJHFK95rUkzLY/W+7XwKPcH3Wr8mIRcsWh3bcArMgzzmUSAJKdL8dAhTJENy
gY0F53G6zdwm0ljkZ2dYDYX1flNEEiwKgNI0xToBtx0GXpCW6KFqwec63JqK47l+
1BAMLr8alkmHO6fBkZvUlzTBiRhQBa7WVhOCCPtUWzD5aAMvQHfYPAs5g4g4aVxk
oTldKhkhZmehGWnJ9OfdUbUziy1ca5/8cXemef/nrJq0XWKQZxcdCl9MaH2ImOEu
tQsRDYKjLZ5AUaZs2eNnde+YMaJS+ptl9nTxUGMFoBiLg5o89oa/cLa3DgXd2lt0
0LjY01mYtQb0VHZq4osHzLJVXBMgPl/O2dh/HEpXfFnjtjJCxTxnTzqX/2V6AnD4
lYRR141IF7kp5FV1Lt5AjtdxlGMwNLt/2bLAbIOAbV8NyIhN/rnJLbUDsSeFiPlB
jOvUXu7/tmDAf3knw9Kyd5lxdFEQRj6Vf1cVgP2JpcJbVMte8KzXTwX92Ruvkm4i
aU+Dqo11zwRB/C/5fS9bE1XOBzYlpxsbhh0wLGe8EN5nJkolHvc8HrJTKI4faF29
DYYpxDJe/enRs08Rr5b2HPaaLjwByOfjLElLjvckYilC2Ubf0qDLjY8j7hcWgUFV
mZTrYwZgLDfeszsSuIBoSLMBLvrWRaZL9NT6c9d4Rddjnsu1vPq5pnyJ6j64wUMR
RzYX8TETXfISTwhak34AFXJB0njkDubAJVZFDpHgwrUW/gB8TgwkSGNKp04xVnRP
omu4mw0lFQ1GF01OAFNpff3hZb/9Vw+jdB8SSN6QUUrRS7YzXkVaBn+I3g6irVni
iLTELUw9g7bD/RMPP0dMCwS6JeB310Qi4uEaNg8OB9WRFJTxG9VEl7oVXweHc2Rj
JhvNvewr3BtsuvRi9+JFVkkf5B+TtrPPTFau07qNLEZusz3mu3xR/V2sfb/4g1jp
i0F0HjS1FD4NWRlsibGQDiUlQtphzcvwsnmchPiwnugj9GlrkxjJ36mvZwvmQe6Y
B3jnOpI2IptPQ4sJPfnUjKCcH7uUqQx+tJZ2R7hesr2t+9YlTd7xLspDwHRci1Vi
/8C/QaD1/yoZtOs7ZYB9UlaN3TdYCRWuNCNCd88xyZiNsK/XEOokn/rWYavSpXC4
m1Cya8xeCpwv8DrZxAbfmJcaL01lMW2e+Ywp1kv3RIVcWdLpxsgejvYqxDqZxrO+
hgydhK7l77vbU02DGnBZLZoroUQogiiRxlsaU7fFhXmfR5c81NXHEJfka/ce+L/g
MInmdzN8zdFZxUeVO6VUwVDuCuKP++BfU/wRWB5kvT8rVSibiXCNEcVuH9RDIoQD
ChPhwo2j+Khx9jY51Rq8H9NuODVF3Kqazcq8TUnpjqLvFz9rcEaqd/Ao7+AhlufG
yKrRgkdzT8y2jgrLxZv31S09do8hyLwHDZlEcqcjlP0n7j+FYc95Ev6a3Zbr6Uqe
iBF4CH2kVrLV4Yga1CaJiye0V1UtmuQ7e3ASpeTdJmytxGs/5/oGQMj74rxoiG7Z
3qwt8YHXtsfLWu1hX1AojzXhFXaVsHXSs+NOB5QMvR4wvLL8s9BhN/0kIJroTCAS
U4X8e8diEfCvIWbfrp3B2770lnAPY0fOfqiiiGIlpTuqSWaalmomNhf5ItHE4rur
5uRRYFPMqkrbygV4TpEL6v6cOJwB6QIBXr9AocQc3R2aEvaN8Hyk6CFfSjSl4u6a
2gN3VHlE5bohir/livbljmPDVSCWE3l1hLALm1dvErquhqsgYneSNNvv8QGPrXp7
tqVIaOkmmg6JtaImKMN0iu3Q8ah9f7TMuEBaU+XiBlMDXDIf7hDHkJDzJW0/V/lM
vQ72u1Sbk9O+TrAeXgI0DO/yjbslRjwXrRAmNaAdDtYZDesO6/dXG3QDVuOO3i3I
feaTDknpoC9UTyc2SpecJQ9mFoDY41ISveLC3rpvRXwOVQjjGJAQ9ZHJJfk8Vyfr
w/PrJDIZf/6s7KVCBGbkdeyCMyCBkYj5OxecGIScDgTDjcTuSrugaarTIF8P2uHu
`protect END_PROTECTED
