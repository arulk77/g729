`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD3m8j9bUc4ieUGplBTnvcw4GZFk/80WmphuQMhoQR3R
eS3m5UKxmcvHAMfFYxY8ou/0YwbHDIZG7hI9rsFjR+80i3K7RLkU7h5D9ZqqCtoF
gws6XgBw+dFZ8Lm6qyhqPBT4QAGlc4q8pGZXZNUpk0jC0Dv/UyomeY4xPQ8vX0de
`protect END_PROTECTED
