`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MuJVtiO1yUXNixVHgaSJ8OscvrrXExxSzBgjWlvppS20meIrMtdfnxXm0pPnJQTV
p7GOsPamWJi1VpqPLoDLsy7y/h7PZsxHGnclUohP18baIUT5peJscjumA6K4RBdW
Xn5fL09nDJobda3h+OPkaGVr/2Joz/9peXqXapogYUb9CnbZ+NPeOpbDBelF6Xv0
lvolc4Q37KYDBgb1Avyc35cWha6dsiKnk4Lk10Pp43KnsDAqN9smAnPIJgsHeBhP
JeAR9MN0dT+03eeMACVDBoXMNNkGH5XMrpgf0yms1D94dTLziWfhFxYvB564w45G
SgowIBMnLIWTUJObyyaxrVU4NHFUGBgBE2p12YgdgU8XhAQF3E9wIuualJor/4L8
HRI3gI+Bgra4HUq1Au/sCYBXkGwt9pR6l3VwuBL8F0rkLzxpxXa2gmT3Mi6u9RPC
EKP356SouOrauFfizuJPNqGNdU4HS96zU0XH90K9URPqWc1lb4gXd3A7NS5quk4+
q0kcMljUssKOzhftZ8V0JZRlmvSXPkQoL/Z8pTBLrH2Ew25WK5IKf7rbAZHgSDGt
MbWWEj7Qt+LbEHhqXBjklBdHXewrTikmbAmsnmBfHgnegw+Yb+URe0rXb66UsGwY
32AfT6hejSKzdk1dXrUcKlKyN1EObGMR1+gJ51gIVE2OLNwiYiKsZLY0HJPX2LNO
7ixRDfXxkGV7nz3k8y9wQA==
`protect END_PROTECTED
