`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM1E3Ozg+KwuVPx8v61g6MZU+ApuPt08M7UCyqksBSVi
FiVgR1a77cgspCXveHaNOthBxzyVqyQx51rv0O/NtVJ+RQA1R2Dsb1rVQbEt/+Ue
5EagbDZYKMNI6ubhnxJ5IdTQFSPB5lX5M286T77JwV5BomhJ9lmxS5J/JH3gxuJS
kmQIeMngRliiosmOeFUp0RujqLSyFZtXOwC5vI7TdCqVjFzt4yqyIqLwUWzZarsC
Jk1mW5yMqXYhWXZdig/q5XFHPoSWNcIR3VXbGUegtpM0QIJ7QYHM9UkoGUtpEWzc
Zo/iLsfisE1pJTYYtMDB5749kOUmyCZ8mm2k/WDgOyi1zz6lsSe5CHMkGUVAzhLH
kwOYoD80tWNdHEWbqwUjaHk1x6L5ym+9yMwAliy5BwRjek0pP60LyBrSt+NzL1eQ
QLwN89Jie/rtshjmF6wFUTuxLQGRic4ABZOncBl4I3NnVLWQPsE1YdsJRiZ8cl5s
k9Sajx863ggP7rNX0GK638udskmD2ep43NLBasl3hAPRi/4eezS1Yxkqh3JeJcE0
nqfeRLi8IGPwsUIQHqbqE3sd5QiR0cFRUX+gZs/49on87qLr1DsJaL9caue/sfOW
ePLeNMZQYgYyriYA4Yh78qChICu98GZambmiWmhSWhYzc7OgJB5uR02uJMr4lBlK
+kAIHqf/NCKNIkSa4it5XugBWOfoCWybmUJLfZdQLKjslRaSy5yR4IrRTBMRAKa5
t7WUMetEyxVoE+Yq6ZsNq3+rz/ukXHDU9IeStI9hiRLX+dSIX1fFTk/BfktEfQis
qMiSW51PL1CkBOBeIm6WegK2IpSpQWJjduFh4fLRp58=
`protect END_PROTECTED
