`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47JSG3kteUpjsIsfAnytIY6cUasi/yyGZk1XwxTg/OUN
+Hncba3jbv9bX+5lA1R6+rW5xKkH5r5NjkY/HiMCzbo+zqJVUi3Sj2HXdER2ImvB
9S/rNOmiNartMN64s4+cbse0XVZmXRqa02rPLqBooNRmQvaE8evQVHZ8Zyf1bgb8
k9ZHYp0baPnpHqROAooh3K9oM5CW3+m8aZsyDv5rqK4uGHWwERkN21dypz6LYLX5
e69+AIxU8bvhLr4hslM+GtlWXeZffxPweMi7EwBfBT1Iw7CZEfJ0hss6YWYG5zsI
gW1QCXYVsseWh+gvbfFQzkTPAEifxyV658LksBeip9lCePNqRenWqUydeJp0PY7S
C0RBEVSldu2QdLkABJx9t4BA9lNaCFZPwEu6D31JbeSlRHUP4YSVU8pCE4MZciJr
gn67E84NUgDWnlH4kKCwKt/vdQOpzd5kJLsmRx5f8uyddzYEblyFlcbsWTHhXbEc
hrSv44W6P4tPTZhiQ+gpHV3EKt7IawnP8W2gitJPk0x505YSLl6dr+IeM0HVMdkt
RpkvV9upJMupHcxK6Ss7XFyY1DR96RdsMi9IfIyjWJ4zatfZe7n18h5QTLB4kYaz
`protect END_PROTECTED
