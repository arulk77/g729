`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aaWvGJUrmbV/X4esVTTGpxC8dghxoko0bsrgLZ/EVUxE
0F+8NpUxQub/lRNi2sB8vkawcyaU//KP8Yc897CJ3vaXocTjP7dZcHZFk2wiOYaJ
0/5vjKJkpk9fP+AlO5f9WYb8yBqq6ORJUc/IMAK93Gt4IUUStim1ltM10kHeTaDb
hWv2iWDygVgk9HPtAsCSosw7fOC5KdopWhjRnsbrxeXe7IKQGcy3Uh4vIDZgjVl6
zVkzcqmlbEA/GRDfSdQEGG2SHSsXoHcnjJDUHP1qe8BEvaDLGj/EMt9SKUPJGcSO
7Vhpbm3BmdsSSe87yNxd5y9Y6+dZjas2feCdimvJwo77NWIS3y3/hX6RIHkHirsx
2d52amYodnHYrGQrmi5vaJpQ0oVd9+UwM70OPt1k5Xj3YlT/CiH43txNXnjBs2lP
x3Ldts92Y99lvwpZhEy1TI+44bZiPMsUJ3bPV+bSZRQvC0h7SiOaof3nTslbWJVp
ErRWCO5HmkLDyXJnnRgExYYL3+Z4Pa+UBFQGsEC/TigcYhumm9dF4UTOkMNzxAzm
0ZwuUWyS+pcK8OTMB/FbNdYK2mW1H4oXPX/pmyRyUl/+dLeS4FSwHClkJrTGzJOi
DCLHmcHcfA9mcKEzeltjEFwj1vdtRQmaJf13Prnf3narWjY0zxzZbAKwWs1TPNB0
67Tr6jWUlJTF1U6n0/EOF8HwJAEuwyIOOI6wFAGZn6Pb9jxNbsKI7hf6CYNMCUpB
cv1HBsCdWmegMRnhgfAp+QyIPB1RW2HVR8SMBcI1KFLpMJKo0TlZwTLYZff47y7H
GeZT/bTqbZWbIYWyDZyZBp0Dik2xTh0TUkWWjB92cMt4cSRLchv32+IfleipCEWu
dm1e+7pMqHJkiCMmDNFi2Bo43eTQcJCyikE2wlyXmQqnLeD+7dufBgI+6NxXOG1l
/OY1SAFtSzaX6V2er5twx+RT/XCF/p2EarjvME03Q9SfFoIxI7pJgfAFgTs3q0PN
ryNFHmb/vKi7ys72oe/DMQD0mY6ecc5h2FPPEpEuT+Wb+K477Al/ZvdPis4fAskx
Ru2xLGoLb7IMciLpfwAIMuESNm7DVovIlHjx/SwDiJS3lI+3JXono/ygA0mIl7Yj
F4VqvBRi4DODGS+8bHGwSB2pLJ9Pyst28FeMKTeDOcemelGNqpqkqB2eXYUQbkho
AyUwYxyfRSKEd4n2TOk0/RDL6A6aIWRx4UV+1HfhPbMOX3hoEeO13RrnvQf/Z/RD
Y4eyCR5Q9LgzDNEHwSfpsYYJ1xXX4y5PK8r9c4dAzapoIPXH9/coQkkWaeAou8G5
GKpVYdELxTooj8jd4w8ZxC8JWbpPbPqLZPDfjWX86TDIgCZNw61T9ZhXHPmopC8O
GFpNQW9R6HI0sRHCl/eDiEe3SHU069dWbT6fTRv9yzKA4Dl4ifiHD2TjnSVjnYex
8I6k2up/bVyBW1oigoKPj1xqgB75cmRWqVLJ0Hc+wkkc3Pfqrp98ZX4aKyPiSXFz
bFdHd9LV27ttWxY0kCPn6EHbAMkJF4hyATLOs4JWzdsYEQoMilmn8uexEGMqIAHN
OzvNwoQPL/K47ZSIEd9FVj8Uj1CBcZb3UTUlaVchNXUUjq3oXwMHdQAZaHlHJ64y
7fk+kRhhdD+zKtGczpa9qhr6HgWHiXyV+EPGlAN1CqZccXlTEeVYHt1jg4UP64uF
hwTEFvg756IWnnV7bwKmPE/WLXe/YBfzlAMZYDZaxjBai+8p5ncWkG9JsXa+B6Eq
2MB2aT2L1t/Q5p717gf961ABZcIfn3FTLU5X6YkXoIpXVu7z8RmWAwWwX7W/fCTI
S7psFiB2EXs2H5VVnZRb5RcYUm6+Dh6A4/zsVky96CP9FvVYTNnpjgpdQ7lCtjSQ
exfrCPmzT2q8hwp4g0TaFoDmFGR1ttrrNV7c8SOpVLDYB7vmSjUXzpHDYP5mGV4m
wUiApAyOsY2b5n1j7thk5VWC6UIyky+0SDBQmxjn7SGte5qMJH3gbjmpjnpgbAY+
Mz6nDJ/PZm45gMA7YpIXt6qGpbNKM8hQ5ssG8e3RwSCgHfuBD4tOnD8IWSJ90ELE
UsYxgUU0DGKf6KxYyskbck+/vEFWf81veT1hk+Wta0lOtpCmIzxWlqYZcdgSLtRv
xLkFPa0eBE4jkSpk/s3XXVirv+9+eQBacg4A+LbF1+DI4qVzXen89KC3mRH5En/K
/orc8mK8/KVHNmbA/svIq0ygq8E+7PSS6RUGYbH0Z9Bpkk19gav7uhIJZEflUEoE
MGGFWWnhhJTGh9MB1E0DMZyvyTHMxPKUwaAW4dEaQUAbRAfkytCpfkNFjveTR9yj
mNFx8gTe21Ywcc/so1TkMh9UsQFO0ALqiEWwge8jnBqYA1lqiN1KHjgOwPN42THG
mQl4zHE6z/W64eA5p3wmQuO8p/cctafd7e75NsAB8IooyhLBoZavn0WofiWXUToD
/uTCIm8IOwCD0Ont6S8HGog+R14GJV8Np23Dq8EvCw7APlEuP7bS25bOiyZh6jHq
Ui2pJRZiApfuGu1ZuA/fsM8l7an/wNK7rVZbXi3yqxBmhCzbm8NoSZiS5mCGuIhh
XXoMG5gRW8oBh8TgU3HmqVHCHdZXs25JhlVP2G1qzvJE4K5jWnw4we1FrWpk5+c9
iH4IEV2//5AkbS1SLQlrQt5Acemytz46N1pU8W2YVdj+H53o2xFc17Yq11pQMGhQ
ByYRJK4LSFGkXZxUAJVL2YHqYT3EfiIxgSxM/6GrRVZuX8lgOy7dK6JQvwcnYDqa
RrEtUTm/BFGXJ98yuYevCGGNR6UH87AlOpyXGprPGu6fkrhHKIDO6w1N6Wu8MOSq
tlfdJ03IXJuthBb5ae1wHnfX4Wc+OWx74iFAX6VHUp8K4cykAYdS25NSA0SX9tgb
UPqfnt0aryYlufkHvNY4iBzdCq99OeBhqMTAAQbmXh23zkx5fir1XzRkskt9YhSY
UNETreCFhSZhmFlvdw7q0wM7raYSYBcjarXmOBQb6AZMw06zNR+yPGS2aVIJD8iA
HD02NjUWEow2J2QwC/1uX6Qkrh2NKI5xrDkpRorfcPv9rLKURC3RJ1A88aDN0LpG
waxbD2JsouhB59KlIb+Dh6toaI0y+9lUTu3fteOIUrwySEbqtzXaOqqDkHBG0IgX
8aeq9MbjTOVNxeI2Y9wUrMWGk47e5qcRoMtJI6rbhmQM/VaT99SGn1sxAv+s1Z5E
B0qwyeFmn12kWYADp+gs4rvpyyC0Jt/Nxz2sQHZalylbIR/vIKl7IDYbTLvSz5rA
KQezJ633z0JdHSMe2KrEvtnpYzFR01sDcV2haWDzydZNfQom3cX/ql3055m8uokc
JqtFAsHEdCsuRpFfC/090mVjIA7PexAgXAiUfsTsKf8F8ZoSLlaVbC3tRK6Mn9Gt
gYyUzVd57ACa9+F+XKWquo2qlX/9sbZpzkHHmLjKW1d1hNrqdMz3D8nprLXxqlBq
rf+zXnEdMn+YfjMb08x3dYMKHf8M8/Alk/VFyCoXGrBJUYOdunnemDtRpTEMR6jI
y2144r/tDTcr/Q0EbwxYhw==
`protect END_PROTECTED
