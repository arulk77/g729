`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDetldDKghCWwP1gS6FlFlgj7/W1IS7O2f7Dy433T5MB
tJpH/xmc8wwcu0cYqkcuT1akYQnMYQxie7uMw8HcQMZiMgXrXBiiPV7m/qxjWpVz
2qH+dWUbd7wzXJ+2CJZT57/SiEOZ22zFfqpNMdPP8VReo1DquwDJVcJyDbd2acj7
QDp2I86yd5oVCRWKr98K4E4rnm2EjBBj8AOOFnnFRDGZJv4aDUm6DmzEqeiKenOu
jNDM7W9IEetRBwRWIJWgy/OaSQbC2r9EvAynpjw/P911W+2fjHM8ASKBE2f3C6DB
Bn++MMHoVc/0zJEk70ss0t9lKLee5GA1Lfv57n2VoogS7gy1fW4HJRwvEhVzQu4q
mTVS6T7tOCBg4OLyca/lawYwZGgDVRgk96QKFbmL0JzuiOxmIovtGI24/A/XcAJ5
KWt1pJr/7l+vNNgpxdsVvyK5TMznNRTLje4O7UjME9eORmCVHJV5zx1dmM0EPRcm
BOK2oaVsnqxrxMNv/HKzNAipRLJ1mft5IbUKKMabaentDsMfViC/Ae+aJPNPtgvN
`protect END_PROTECTED
