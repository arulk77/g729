`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkXfxxzoQ1Szctuc2bBCBxieVpDWpJOk9M4qvOKYgAffm
vYgDd1h3BQtUUOAePj4Pb/NZQjzC+H9OpYChCJrZZtf4i06QSq9QVG6wxo3glLVb
YaJK7kWyTMFYDDC+SBIl33G5XDcPOBqlBLXZkisrls3yIx1ATCuvKgyWmBDuF9Av
nk6kHM2oIMWLjXjvymztfKGtJf2V5l5D8zAfrz9gduyLTtxgVzbU9TJCk9Grln7W
Bl5G1XyC4H1nvSwxVCx3+B1CmCNB4MxOWLaVLpkyJxQi7e6QTMlt4cKpR2vTSs0m
E3OoMBmiPL6jNdwZ2SzlgMnYk54AJuJAdso/p6kVSk+l7mR5TgGzFRZO4LDBvuq+
hpqk9+UW+URj0e23ZGblj4x9W/Y3P0jH2drNw9mFaAiitKCY+QyXYvbV3dq/CdWO
ReEHKrobYMZV60mqVUKs3eX6Xx5RIyfX0qz3CHs6Ev6B/LXFg2tUbp1cs1MaA2RO
geCwsWw1odwJUyoPIfaf3pTIsRNz3hWQ95IIK8Gas4OEZfiiy3ZzsOZJHnVy5rip
0BCXo/93uSnBatQyjSLSrGaimSHJ9/1t2BSOmGfh683h9bHVIvYipX5nFgFfDVPj
7mq5wkph84bCZAt2lhvZyQlhAIF2T3m7nY2oGRejaU/+Kg4vpCgc5NyI/jSxofmD
LIXhxFvKdJbjPyIhT+m+O2SCbYaZ6PqqpKM671N42UAkbPehzxadwlQgltVFcfGO
Gqrejb3v/V5NQmZ/na0TWRcEz407USYC+dGO4YXN7aaoNHRq3vMZxqQ+DsKRk+pY
AY9BSc0Ug5d8dsN/QJ3vZsnd6bWBiWENSYpx+TDd3kadi9Ya4SDXsfGjR7sXX/gA
cvboRjssrIlo8MoTz2ko8Axlv8L1kVpBHSu8yJyyb2kGg5wTtz3uAZQR8zsR9YRO
N9LmZ94EWF+LVi3GQjMH6edGrdSg3Tk8HxvgIhOaaqRbGgS6xoQC+XMmzMrY6Qh6
DQp81RvRBvGmnM/6a7Ig1UPfhdBM9Y0i+Zu5l16dv7CYainEv4CDWTkwkAswanXb
PxDHDHRsHVe8pxiEEPlYQlY71z/NhW7PFisWOFDzXKM66khnc5gG0SsJn0abZsrX
FbQO8HTUNpqY1R/zGi+3rsVnaycvi2TBiZAInQqdo37DDiGFUuQJ6hOH1yVB8crx
RPsQPMu6lYr4DR0moQ5iH7j/cc6k2MyDk1NSfrj7OP3hrrmdjkTpoD5HHoKh9WQL
iZsgU5PTokJHV54UgMSrIF/Ypa0t4nYhONiNRJsdDTmDHs+MVu2RDmV/LkihCsZ4
SnLHlcUBeHxkxp1w7CjItoxwQbUj/rdFJ40/p2xFHtI=
`protect END_PROTECTED
