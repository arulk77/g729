`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+I+8SIkmzRJru9FzXQLAsbji7ZJdkP5tOnCM5mxfF7s
/qJlFZLeCyjA7Tw38DrX8kUEF+U7D0dXzPHXUWfHlE3JAJsS+F5DGautNjYV916k
TfUM7/B5nqVpy00Pog3or9zN0XdVxXaKO+E7xHXqjnoIMB1TT96V5SaSqLD7Xqah
DvOLBU9Tkt5RTIQ/antnF6U2lHbMtJqLvP4Q4Z3BnHodLJJ+CEFC5ZhGnTKUqT/H
4iDfeYJcFwxsoE+XvGZol3oDOjed32eB6h6okQoF1amBkOue6XICU6D6tZqP8bs/
/boeMk/vAorHB0SKC1gAEIfLPuwikE7v6YOucb32vsfM5HJFjZpLCWYIjhlFr1l+
MXH9qdm5zr8yIw99oIoYtw==
`protect END_PROTECTED
