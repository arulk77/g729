`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOdwybVes2djAoOGuqnvg/9hyMsV44EFXRDDxzsElZII
dWr1GyvPfQP/dZyfLkqGIyXJ9ELh9Sr2+TjZovp/h0EU7OhtFjfT+gChpWd36/aE
UUNyzy7/zVy6HWJIOhhkoCRZ7N0Ee1FQxQfqF1fgmZROec1ulRTkr/BKSeKX28i3
`protect END_PROTECTED
