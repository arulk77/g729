`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG/nkVmrIfnbk1+Ou2jL3/Y6BtSCplDyGgCE5TThE+Hw
pGqgKToYTauD+UQq3e5xdLkN1szmxRhAD8CiRSWjLs1VgWfpCQxFl35BX9/tSN0R
fQZrL5Pqvx+WOTjx7AkSnpVwS6IWgISGtdniiO1xd6yTdILfLBW+9Y3YOplFbs//
j/OpYOyQ9PK+Bv32FK3Hi0nnPYD/eSCC8omXrP+kokLrAgLYOr4a0pslq0qsvSXk
7n0bHHWEMGiVGOjNfzzuEH3Nfymb520+ZAEUqHsMrV0g4eBx5tx7FCyk7kagHn3y
genZL+xJjJPXH5n88w2SJg==
`protect END_PROTECTED
