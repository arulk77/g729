`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFxCpl85taRC3MWCcPrPf7d/GP6Aavu8RXgXAeiaC7+a
Wf0hqt2wSqCs7Thbn21ZBZZolo5N/gfAy9cMNiiV96zkKrejF2aRk7GIfaeInR1N
o0tqjOAEvDCtVF146KxqrmcVWKxmgzFc1P7LMeKsoplDC5zz0Q5DfptAy/R4nVwS
btVUEBzMdb/LXUve5pGa/tTo/60Icyf0BcZlctvuEwapCV897xvQo/Y6aFtLRWwf
ikc8fAJHbKryO7rBdy6/7bKmB5478YpxWSp2Lrks7/pNwWbAiF9SYAjHZ2wb4YQe
oiEs6LKgRUspiIjFo5/cncQQVm1j908LavnfDIsKfzxmAPDsAh+wfmgpFqrYhRAj
hK/Bvcd2oS7fyAauZLJz6mj9InE0rKmVbVmNrMkVQXXlrBoEl+yRjX9BHSy1Uf5P
wOuUWQdviO/vALADeXrrurwbWWJVazNcbnhDI+BVLf5g2Gr4fy0tkYJU+cNQFh+Q
A7FaYjRrd5zXQx0JWceXwSBCsfQXKRffxnVyOigWBnv//RND8WB54XYWqmHRzlQr
4nO7FDTe56fBF6bIijh6CQ==
`protect END_PROTECTED
