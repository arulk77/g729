`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bpH45Z3n30C5YyzY6x0AhPD3pFuc1/J6U2xQTh8gpU2FQYs/eNYKJg9qS1XHoQKM
AuRaHUJt/f5r66kHYBSbR3k+UtGuefrlKTpFz715asv1HfsGkVuZN1KUG0HH2QDS
25flDAuMMATrBhMLwo8nTyFwZVCVb9KJTT8jwFNEu+DgSpcJsuV38zk9YNyWY7Hn
CpNMITzQzV7Esx8CkbsJGV0rtgr1czHpkcS+pQBtAfjmxwiXxiB8Y8Zu4NieUTZk
sfovb/pCCghDUJhm6/x2bEvInOnM1rA8Zv8y6erJ0ZYCe/VfjJp2FV1juNdEWJem
BUxS8TQIkep0Dpo5GdTg34LkHHFozCQWuMeQG17CiuPAaVXZRqmGMmkeOWhULf+0
52UbcchvnsBbo3QmIFVaaDkEPxkW2wKVdCwqi7uL2/d0+rd0FFSz9/3wDDiAKbLZ
71988gKJ9OyPY5wEbgZNj0Eb/4RQFWbBXh4Dhzqce6jNwUwzh8kT+li3FPr0xMJy
ikb9qQ+GUWywvRpyWkgyPKJ+Qqz520MuIIK8brZrh2n4eVu/hS9WcApnDmCaTq/T
k6jX0knhSn3+BE2HqYHGEP7oLukYYXbQ+TkcQIrOosJCroWoRt4HSFtOqo2VZvkc
Ez+dz0ng2kK6+TNQ5y8WSCAKd3+D/gadw8iqj8IzDe1OrTIPl0MTjr4Jp2SwD6I/
7Uz5M9pToto96NyQ6Cw1BcmpBRa2BMqgmd1Fo/7VBqlcjOGyhM+g8Z9QJhg715yl
ErCdDMz343JHmIc0M0NHPw==
`protect END_PROTECTED
