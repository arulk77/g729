`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBGdvMyM9eE9OK9B/CI+q18/nryOv+P8gisufD3ssPBs
GIVyiMPnS8oH4ztviYrJYFjvgS90Sj2M1hetX8GtHCXri7267a2O/AGig+HrVldz
pXPBCHXzwhm+nOAybBKo3BwvoeIRzy0OAFccZ71VMvs/VnHVQIBAQLpXCXrEtSPP
l1qlNj8PJBViC2/48xxYxKk/ospTd2d2Dk3xJUPZoqI1cNjlQD4v4Vlycn0p8ozK
NAalF2b+cqxj6hIx7q+smWF4LXs/8hg7pUJbiEkQrXf+Y1taKqE2Q0j2o8JQwDef
KjZLtIaqIe0JB9+lF7WJNJzzXwFsML9rFo918VJML4PiQVyv99tTLulDCEFnWauS
WvFGyS3VU62MAEWDHPhszukuLKzirHKx68uSq4bcodDSDC53v6jE7pcfwrR6Yb1u
y8P9QJTvzqvsI6GXy6+sr2LXSYCNu+OIeufTimbqHOPND/H7/m2X+QcANRU0DW+w
a2dOn7C/A8iQF2vWOR1hg+9/tr70di05jJTcn6DAEMSAB4khzjsEWFOtJVEMQVP6
`protect END_PROTECTED
