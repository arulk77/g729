`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJdGvMvtnpZNh2EROMOMDEyaJrmIGesr8ULTY25FdQCX
XyeHNZ66393+71SS27gFHm8JRt4EQMe7Jyn8TWSP14XleumkUPYV6tPS15AyRJcu
tjWkBv79bLIfRCFIp5Hu44qhi7lEXVvaV/FS+fINXAsKFJ5pWk4oh2iyCkSi7qgO
WDeoQS+b/SKJi7L1JCQ/0w==
`protect END_PROTECTED
