`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu433pSsIYrGd2rl4EBniGG2ubFO1jnXJFHrhfCZzl0QRi
lpWOd4GY5avD2YrMb9/VXcATy8TQghpR/4s021tNp7Cb9F3R2KtFFrrlxxxS3jeF
KtR47wihMoDiCJm/9OnA7Xagsyqgy1JMHDkwqDyBHGvzaoA/sO6mdXS7lGXzourD
nUR6iT7xzs0FzgPXcw/fgpZfSWFm7fhcpOsGFedH8FxMo3SdkK7+eKVhGFNcO12V
QEVssvMGSw4zvKK0bPi1WpjenP5BcTt/oJwNb5LABEvXo9dGXh3bJ1o7D/LzzYP1
fKpCQ78TAy/diXxpooKaoWd/PRfvEAiwh6R61V6mFtDjx1SVY3plj/KAAfGu8oyB
1KUsgi9W99uDS5h13pRyNw==
`protect END_PROTECTED
