`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO7WUNUl94sCVjzlHljXoZuNsaWAKadIuInVWA7IKQYv
SYEIpfyWzO4VikpXKjgCyEnKyDBug7EhhFKxHuew+GtJ520j83s2ANjboDa+z2MB
Px/+ZoFnIiQMZlGNT5w5xLAZlT8ZkuS4KuLdxOE7k9Jip8cVwwjve+W96NYly5KS
M+1Ox0dqUbXCIw9TPvhsizVmiRtXS3EBUe2UN2FYmlJtpoDnbzYBDKSBmMhM0ooF
jNMEYjrtLSm8MT51mT4vZEXPq1cj7j17vUEYI+qXFr5kT5ujEIcVWREfxOSK3lkr
wZ1E8dkf95mvANTOTa8Vfg==
`protect END_PROTECTED
