`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN7QnUdSB78ZuMr+0lwHOeZ4wZGGNcygHZSUzLSgAOot/
lCd75J3PAp/gyImerV8HXGZ/TTdTzUSyd/9PApLzizZsgwpubyxqNWrsse2Ywrvv
fBhM7z9SdHR0wi9t3hfg2iJ1dgT2mqlPevzYG7ttOZaRJNPfMR2z1iDBRmcUmoSi
lQukxAIJYYrXt6/038QWg3Jd1pql69Jy/vHpYZHQeREQOZDzQZbhcZZoahEQ8bi9
YVugdEzUP+PzHtJqDF1Ifl5zksN8T+ZxkmaRd+xiTErdqJ7X9rjpreH0s19DKi3s
Tdrg6goeHDlKkYCAIBEVtG3xlM5g/n1MVXDSMu4bBKRa4Us5ioM3OR3AroysUB19
d8zTQv2eUMiPiP/RKch+CHkbfYs6dj7D8L9LJJpNW0Vl/QworfHzBJDu/YYBPpBY
QBC07vuhhbuQvZv7BGI1jtaXe0lcW9DRHUwYc7tB3lN5Ea56GNXF48/ITdyS7l/9
dl1/wW31Y1DHvjRUGLN+BLW3Yy+/GTvWnGevwuudL+rREf4tpLVJNLyWjv/ONd6I
QDoVl1C+ugfZsP0lZTp+8ROIhbM2TYSah54i5LqBEbE3R5KwoxEYhHlZBleyoQ21
tEFVmNZNlbpizkVupiDQ7xiBJsDbY3ssE/bV5s3Ro3Dz5QKb58PeWm8NjlsYh9t1
OxyTPl/Yqt2UbIthQ9+sGTLKSx9DVFsidjwx4q42+REqq/pZvYslfDO1Jblq5Zig
oKMJD1BPqeMslTS7aRxisw16zlfmm56OhlpL2opM3j5R6UGSxT6n8oZnv+0gcnBm
P0SA9LfWzQl8sIcGMZ1VV+CATJzUSjB2n+Pbzrlk8NnNC7F2D+K1XerCJ+RmNcxq
yWULSXe98uyCVQk2psweJIwaBlDqEERH7iVyffE0B22h5UOEPFwrZT2nWKiOV4o8
63PdGaC6CSdnvxZ9QBvB6t9vXAfZxbDKEMXOvOXud+wY774CCM6rpk48Y5sIz5BN
3MhAx/dnpBq06P2+0QXPSya2QWFL0EStJo4L9nfzeu1IhLkxomho2vdTlGGFepgZ
F6/IdFBhG54PQFzQdqFlLhW50o9SMkOVnaT90jY2gfwypoqEddBg1gu0+8zO1yYE
esxuiFOKRtp+0a5LHbtDX2DEJdrHKeWlrBxS520OR5miK0kwvKmuk09AQ6jcMIee
QSNMAhC4Dm3OZoYWxL1SIIB72WXCR/56W/F4OkhGd4nqcCp9dlEB1pJpYZNuLc99
biwYl4zpvoB5Gwi/gmh/C5QpeoPYwayqrky4WCDxO6WeccH1Cwl5qDHx91lq1i77
18lRPivCPzWnSIoMsV03ri798IDhZOngAgGf7mSFiU641KGxzn8zW3Pl3dkRT2sx
qiEniacYlAwpkV/8He1FZ1gHBBNt4XTg7/BwV1xNsx8Q0V+UBi4lFxk/VT4XnbSa
pw0OKtZNMq4xbQ17KIIkuEe+ZA6awk8fw+IDhCUyzLah3xtFA6LKLXZsa/ylJ9Bg
ejjPCYoGLr/05AqIULc3U6/wJHYPicnP/dzxupSVtZb/Amr7Y9oR1rayUBW/LtN4
phJnjQHatcxlWvg0UoiyGISZ+wlMuym4zmDZbkVJLTNeKiHnTdkkrRiObTvRS+v6
W6r28eShqb42eVyLGRnafWZK8zUO4eWF0RvxEZ13SqOZ59fEAZEsroU2RsJaJwgT
pVlbEYdui8Vq7kvG5RSInVsP4UmyY+K5omqtc7+AMhbob73FZYfW57TCj/DENjSM
uPpRKaOxSIVipYzOUoZJrwUHWmaXc9XFMaD9SrX/jcjsDNgva1JW0Ae+AN/zc73w
FrHw0e4j6KR0OIbd9sJwo2nkk8TFxya6GIveHOwtB9QT8z3dzBBw1YunlavzeKKd
QTXM9610FH0Km1RCQ6hOgS9wAg6NlbNJMS55RFFP4jWzUZB1kUCWAEhJcAyJ7jPP
a8TtvcJ03TuIYuukbhde+lSVd5RdHamkCKy86mLiV2W2N7dJW6y2/odCL1iUpkbi
BM9WCFds+rZxGHRxYpLovEyWCQAPdogvaw0HFf3P7kcWvBXjHI9M9yCsOksEqtgB
2G54qcHulnZPeWrMc89rWAIrT8OmZbifmKN/bnp6XheTkvnLDHSLNRfbL5EV3ySv
WVIR45g82GJHCV30e2L1T5NpMLLpphyOi4GAwQ3QRqi5CVMiwsbuAqEG5qJGLx8V
jfcVBF06M+aijnNJqYoJCpLFHELxJUEoEecsE4/1DAQEQzEcUpdTaiEJ/GqoOmb+
xL6RLsvB7bRaJ0GLnBXtCdX+7FQ1JVUHZpekBj+lbeme9A7fuLwCVePjhC8HJhk6
4hGs1cS0+iUqm5D/WwlRxGrPb2HZNmm403BXKlqV8qbMhlg3Ir9xiKpTvnVSDf8B
SyzTmjqYn8QrXiLhpLfBohOqyUdhFRaRIDRsngW3LnLk5E0OxnKj6lko5A3vGYEd
HAbg2ZD4ACpdpfG9AjgTBiamyCLkGpP5PxU8L6Gg3PcJTWvyiX78Z28BY3jMphm/
G9s9iVvqGnbeRO7ao0yILJgd1Kx72a28c0fKhYFcbmU3Z6UZMpbVyI9x+lM9CpvU
f3MR3YE/hMsvINu5BbUSgg+hifHxGo1q+3y3t6iukPlPVWoiai55mH8C8hMaGw37
VjD7L3yZXSA0C4Vu5KcQauIgRSMVvFHNPYUO4Of/UX4E0aMIqDABHi6vUiM7UB4K
IvPXOsukasTC1+jQ2PSnmkRU2fQXMSmqf5ST8whOmZAdgBwlXHCuN3SDBeRjpCA+
Z9pJuY3BQAUkcvrKht6iXdwXxTjwX31NS8yWMWbl3YhQabUvjAEze3c4mHjwG/wW
b95Nz2HIjEmn3th6tXxVkBRNGoFtfhdTyth1lHZwvGpEF0CwxWgCWsMGqrd7VEfN
B8nVhryVgObwBhR8IthODFrlCsakoQ46qmvb4QBy7yJjuC/6W/IUILp9uPMtEt7W
UD6RvudMMY7CGNtQtEI5wg8/QcoeXE00zaXv1r1znoP+OFkvb9idKfJvtYjSXX/V
mQeerXFKnKm97wkrW1WhK6teey8qMDuGEXzZshz7Dy2Er879rYqOA8dBvUYlZMis
Uay616pk9S75hkk5vCw2KTe6u2eK/qXBr+gx6iECOOpw/MThoQl42pf7CGLexmMK
exkJqKYfpQ0+53bFF+eRqFWmQnTZ9dXxYV6dyp4VjDBCaZnK4SLKRnkWHc8gMgYh
QnJCtCj1v4v1tbbRJbt+XODEyRfYN0+r1NNJBBmfV6DXxEL6jEdTzzxZafQvU6qE
pgHNOfAQ7hIYq3UlgasgLYKph5zDXThgGZDnKrQayshGiGkGp9DTLwhNwvKxN0vC
wk2qJ/CGgzlH1s4nmc3qXNiBIFmJa7ezNNcauQyABSnTbNhtvj42FYg3334GlPpf
IcTyKE5vknExBcpt90kQR7Qz/BlHZ/CzTXNG3QuAqmvwvxu4n9VP35tlzwgyOiS7
CfR++4NM3G/lpCSfWLIT/uV1V57Y2ryBv7ow5qMQkgysutRRh/OSB9HKX3Kexxvu
Ph5GkBUUsWuh4BDY+TJm4VUEsUR/Ym+gBqI7JJmPl6Qdko/R4gLAw3e//LS/o+5E
Hj9H6XFfI38bMjKdCGLNJgVdI/bNibNX6++sxUwP0KdNLWxVpXAhvkTbFbO6loHw
/CBwhVOAjozGb5/sG+SNFU44GzGddNn0U3DnJqrtM0fsuIRuE3rml5JwllqnuCa0
lo+xNxD+i8QpnghKrEXp963OPrhXoCa9WKhwmkDkiaUS3mBDF5VP/ClmBS/2EqTB
YvhBGEt1HLxFUEOOEIRJ5adNO12JC22nSPRZMexSSvTyNj9dGGLlkh0icTR/on3n
FAQP1VNwhRX1kaaeOiOJBzmrB5z8GgpS9i2B0ZIL4UrdWid8vlCvwPkf31rIyxLp
MXISz6VoiIgPryTFVHvM1tzKT43Mdp9aiDTaoV0YPCwKldvh1+mQuTvqHR1ye03Z
SmPcjjFbiJtNY7SJODi8VsmZD9T6xpX8+J95e9jPEkBIc9cx3waT/RFDD9P80mbs
yRE55yO0Z44PqOVtjqEEKElt22FeVdFvO2CKyPIAZYBoOfX5RmCm250wJAvINla5
K0oDk41eI63bwY1sBLnKLhhdPsujCFHYFJmwEZ57EcSXyxU82EyXXbuhbloJrMpW
EhMdy0fzk4i8IrifOfn1eCKXyxEYkR9XQnMQQm/8I8aRDKnH8+ZHw+UCRRgj0J+A
cwRnekeQCzhQ2gQFV9V9SY6SZh4XccXqPeOobHldsPiRFLhOoo5QWZlu3Flc+GWP
ZcuuRACa8ncsPRLhBCgJfV18h5wCHMf7KGFQIHZwT+g=
`protect END_PROTECTED
