`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHfWxoBNXO5QWywZa8MhRJJB+DMMz0p1l3J83iR78C2G
UO9nT3cN6P+EbRH9NRTN6xOouAuuT+ttjhdVkr7AuZc4xbpOl551DlvdzbR/TWUi
pKwAraYH2PmjDnA8fM71SfgTsMERrZ8ADP+lFS5MSgeEPkey5K3Sh/702FzZ7Jv2
YVjtzjXw+OyK+TeQCZ5RDKxdceIVBzrk/Ou+8htatpZ+cyM/s1L5iR/iGoOozNOv
7HhIHraoyf1qBdma1BintOTRyAMqHqu1tmjEZHcqTM5BtqCbWd1bPTdiSI00iZqn
8aTvDtTODV/7Kdr8hnafeEdisEJJXxrmtc2wwwLn8Zol//XrDOwGZnrJ1jkcX1oU
vEw2FTtIZOb/XLvVn8E1qr9qAJ9rKcwIXj3sBuUxa6WjaLsFGjy7I2f9E0P/ykbe
LuHfTIXqPNLtTzui7HGYjbM6V2Fv3ugprz+m0EV4VpRamXNxi6jD2tH/4w027Bfn
KBTEpddt8OhjllJKYwiD22sy5O3TJA7Y8h+iXVwGRByUv7UmcWVdoNNJLj91qcwB
bv/Uk6hUm28A2Hw+o6xK42bwF78egFfBTPTMZvj+eVrBbTqXRLREjykPSuixoNqC
4mjTYMG1DVxhtNAf6zeguv6iOBC0WyA6ExJPam+4kZfvFvtq/Q8cXKQOmxTajJ09
`protect END_PROTECTED
