`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAwM0q3XFZOka997z1PM9x4WYntqVcKM+xB2HjOC9DEB
++WL60BjTwGvdiiOJQbd48VGvEZptmfBF3b+ucsMCb4SgPiFfcEcY/RqlUAhLVzu
FwOd0eMY9OBgAim3QWE/ZSgwqwuhi4KuQgf1pVN7ODarM00hfqbHEXoAjsXLcmAb
zTKiRoEtUwBAyDShSpMIvsZzg4MmxqQGn5npblfiaw8cJEaN/IHdi+70ttvMCbSg
`protect END_PROTECTED
