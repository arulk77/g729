`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAU9CL9K2MOrG1+Yi6fac9HNmzy1sH4hOzOG9DSnkd1R
hjCViKNSwIggSyxqMD/5Fa2+G2BYqCTF53Pjysjp8k42o29YYVQTQTYty5M83R5E
mTLVxxWR1BEcb0hWneS3AiSPzRTqzaBtnN+kiqdc24m4Op3cWGQiPOs9iiXsb1CB
JgdQqmzQ1jC+qoaz7kblW1N++gL2IJb1unYN/2NzeCss+5zGJlNoedp85Q98Uhuf
EusJBTEZRq1B2gAHZkcEAMs0TuU3pxhY/uucaV+0eE82HKFASwEoDHGfDMi05JUy
6uKKmTAm6OTSziyZjTiyu8VccxGEUGfM7pv2vmYrq1FlM1Tny9twLb3e2aMbbC8C
bCYTiTLCGOj2ZYMVTRCVRj+W3Nt5iVIDxyFclaaO1g38zt/P+mQfRP5ngFQcv/8F
Qo3fyDF3yPWRH/TVg+oKl8AvCYJvtD7LI79IWiS20veFJnzP5CzEk5ul5TvH9jnG
`protect END_PROTECTED
