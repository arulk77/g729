`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN0x7xr/1sj1gWO1nP0d2g6zFRpNle7eS3BCr1O/W2yQ
PFp4DXe5BD2V0LFiEZBVtSzvaWCvdGzicv5i0cuo/cHR7uRlcWUleEM8ftAl+l7+
KLyV5yhLGHIn0w4xx3Q2cY5AFNlXlpne/1I7bJiKfpEawcaoGfF71wyGkGQmf1AT
MzLEswTC1Q3/q+KhO1Hjen0GBe/RnApHUiipSYt0qm3RBQ4Ey2y7Twlszduv2AQj
2OQ1nCzpf+ZzdLxw8T3F9bMbCQGfYe1oZ5za3DPABymPs8flSbkjLZAkuoEKyNMp
+ylN1ANVcBGOwDlhxWJ2meD6/IxmkhQYvZABGj1i3EwFGM+souSYipme9HSE4WI3
t3l/XN2bAD5xb+FCtR7oJFrMu2d0U2JL55Ko8hM13tCsxNiidJkHbLVv4tkK6eg7
`protect END_PROTECTED
