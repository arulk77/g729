`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44F0h1bRAb//OY3dgBbMjnqrtOikvqGiWIJ446Q9XnJu
fEv+eSwwMMitil9KRIyAptqw4U4R/5A9Ri2Rv9XqOA2r6CB4/R8rvDGgSG2n1+I3
gGtonRyGZYJvegbhcv0ZfgnVvLDp/8Z4ockYbZQgKROaPl42h7hKhkhkJmUDdOqa
PhKGTfCmK5d79jHfukTP/TBgR/20UhZ0BnhsZLqFcZNprPtMcnmzSFw19dJxjX3/
4HiLH6H/Qy0EjjhoRwki/9FpHpMa0s7bl2o0gmJN81baRW8/iYulji8YMS/6AoRL
BQSAMVVVKSzKhSsSICcL1g==
`protect END_PROTECTED
