`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAfdN5dHpaEuGLEy/pr73ak28eG419SaS2XTVqzYTb2q3
7Q0Eausl5w8vN4icycbdw/U+SGc/msQmYE49bzLN1R8qdQ2f4lefcF9kxMsQNW0Z
xgT5w0yECrFmb6DR8yFkqSyG57eXqQUipq8eEeVA7pfXyoaPSQ8OiWyWWg/B5tF6
ZElX3hWwPUMH+GIjTehJfGexzTOtYiF3eQvtRh4zPhOLAIgVSdzCGOdkm9hSh8Tk
TqnZommpmxOV29nMZaFMRPoBpit+EO2i/vUlDY2ms9J6ypmF14rdWPUSbqG35j9q
xEGpSKCGD6YYNSHvwhAmz2MNg/XySsTOoYwZmHnbpNUK8p8dm5yFEoePnAVeWETp
h5ch7NyzwE0Dog6yMJLfaDvBeyaeZpKAZovvqQVGQCgRA4Gya2xe2y3+CUskyTK2
8JLO2dMF75O0w+ThLvabZXfIcUIglT4k2ywnUYHmLjkIMxQoNSnB9lJ8RSjRmizq
b/Fty3e3Kn+/ooaEJj+9Bj6D1gdUqQylrllexTpxt6g64QoQsbx+09JZ2YwEB1m4
PZ3mEKBVpJW4q3mDZfx1N0uX0o8GwkFUXtYI+YaWWmN32As/EClIXnlZ0vZqsH88
2zoEG8qfnPPbmIqN1Y9gAbKjl+PM4dsNhwAjZrVhd0IzpPbj9PK/23TxpFwTVIxR
YeXr2A/C3yt3odc2OHi/o4Ade8Y/3SeAkIs2ToFbdJaML670e/ZiUpCQym6jh5Oz
rctCJX/v2jlOMJXW0Azhg3z5gE4UGvqQTmosFajlSErBWPwCiWZ+muns2UlxP4PV
uT6uKBH1bqYy+CFOFJPBaiLrK6LZ2zbbH5hGe3jgQfPzs94U/cUFKBoHBxpClvw0
NmG/iXSq4Ok5ZK7NSa2t+q0MaTpkGRYTzNU15RTKk8YGmJWw40GNbE6q1v91OI9Z
IQourlkaAFM0iQjB/mGMFFR8cuWaOUaDNXnOKEy5MDM2RKrVlEEHBP9dBSG5g2YG
B9AM9mDVuchVb+CptIl0xM8257SfZtfRYm4jEc1WYhKwvATP4BKX0J6UKDAksnhF
Y+01GBvvmRLKamo8dMHE3pzxr6t3SEzdxc4HA4BLqah7dhgBkQh6s0WiyA8cIOrQ
u/NWf8ddYPylgSen2R4YvnStDLB5bcjaFkHPnHSzU1VHyTbby5nmHpCXxALgzylW
gxsUtqNzjt47mRMxKBJEXQ==
`protect END_PROTECTED
