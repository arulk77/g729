`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEPA44EhA2Gdryf3z2XGdYT/Sp5GzHR9h7QW+sMI184a
yWpQ4H/7BbqRS8evpbwZVqCrgH6b8hxekNikpUBmYEsWSC/4QGGAVwNT99H9zp4T
yxlASogtcWoswA2zHcZhZDNI/YenCR3DqjnNLU9vngz8VOgLyPagoVVkkgIzNbHn
YwFb/DZ10jQqhDHmA5CJKNpdpLwlVVN21fFZaufaN5dBsCOgNogIFkz7zXmT3cnI
zzQxuKfF2kfUZWwoFnX1nHXaTxuQhelxTZjH5S3DdfOCtUIYej3ELvyL+7T3RajJ
sRRfFGL0K3GpfSrvHLmRJA==
`protect END_PROTECTED
