`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4dnKHnC4aeN91eoX/NEmNdcHKPZMGq30DyeAd4qctQz0h
WNIWfPYB1ytO88SIvN46aHMaKJfQvpa9V+XwGj4OVwb2Dbkvorxb1ldKf/BnX1P6
rt9vu46sHi39qrJSJBr07NbmjpAK9YsihlPfmzImggzI1J9LnX4H81Hq0SVY/CZp
`protect END_PROTECTED
