`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QdwybognSBMDmJQADBeWXp3ibmYtsffJh1FpePAQztAAdJIrvuY8qoOkh7NWwC4o
suvCoEnJFTX9ddNl0fP/R06HS/CtHwucKZYHFJpRFquHo+xqWGFVHbK1Bgy7LL6Y
IZ1H3nW/ij4x4X/x55rtM8O0S63Dj0Bfo3TAVrRV4XRrG3tmsH9RZD4DDJgCg3EO
s+mHX8GvLE5PYFBaHUgzxfnXBjFC95KrytvGQcjv8iu9qKpylGC2WsfzDx566wL0
cLoghxjnIRSwIeLosAIr4HZ1aryMZn4ic0zY2xkl4OkpoHNRkKtI26BxICnbTXEJ
9TV3JSIe/+J+niLnqkdBrKAhMynGYSg8raWw+gqIzTlEje5aTc+1a1UEtA/k3o3B
goOTrI0zfEFQwfjdZF1iqyvs4DQOaMMLXiWsvRyQmxyXeETXQdiElTY8LnsVxT9d
EDO1O2TRkj6QXElzX6TJ95UUpUaxEemYuTXnGUrLbDUcPhQlgEo+hgjju0b/PywX
fYtNo7UsC1CPAmdsmg5aDGwhOnxFKwPipedF5YnVqS+ZuEyiwB3ETj0LtFQLKLiw
p5Biay6jj3JF7AwoDdEVy5FpQ7PujbsurCSUaHeOv4FMO84Lix49tJj/XEOR/C/E
SfVaHz6F7edcCs+GG+zqgDxHz2UoJEQujMd5kCFSCLpy7LlCYi8bRb+1siDJB5wA
FQdN2urP9jLL6EGOA2Xf4DsRDpt59lxgR2kqPZNFKzs=
`protect END_PROTECTED
