`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkTGsbOmjZKjZJb6/eLY55QbyrCAm58wwT0NdOL7cy4iZ
Ixk0pzVALXaeii4M3LkonGp8HT7w+WeD43YxaeaLiVobCXnV+jqy16nKLAHqVzPe
W6/y3TkseGU87ryU7pgEUjfhO4JOGfrL4XcWqe/wOsDfbyo2ibiGL/dSupsDrF8D
2YTA2wKo+iypreglbfdMszBszRwJWmivfH5x70pAy7D2hSF0nsz/Tx5HY77OIQpo
b10j4yfQ9JnxrzYA4sCI8sm2jo717J3xyv5BYkOtkivQGjCMSgF/cYvowZ/N2SO4
OfEIQHwVA0ih5Zaoc1qm2GoNE6c3+vBm64SvJ+1oZZ8fXDlZHkAfKPFWnIjU+NHM
SkBJPrPIZIjtF9XIx+qDtYQQ7H5MZQGQ0G55galaz8MoCtmb/TtwQB3dQnesYLKQ
4K6P6Oe5aH9VOC6VSOERaGqTP1UQCAM2YzNjuARGtGjBfN+AgBkMxK4FZJ+xum0A
ZBv2kwMCoXMhvJdEWiOSkvZ/3IXariGafA5NzJ25ibP4eUlK732GWvxSS+ktBJDN
zzpgcHNN9G3kiBoiBxrPD6AmXF2slM9mW3BzB5+zQSgK+gSkuc7yuQBL8kBzSAxF
w9Zg5blKnlnwnUu1nZ/P+exEJI44AEROIFVvgdBh/y2uue18iU0synPJTH8TexzW
o1XReFgWgC8JcU3EUqphTirVEfDHRXQvIp+P2tLQqUTjLGO7RgZQAdSS1R46eaA7
woVLHNSCoMXqaLMXEW/r/gpPxtAu80qcjWLYVXX2syIWhRlOmr6RwH3ZL0wUL7xi
KJwqGzSPiPgMz+EmWD0Lrl7NSXQWFi2HfbMsvj2b+jm6k/DpLBoMRu709AAuQSca
IfBCFbCghWlpZCQ5+z5LpUWKHZkEElK0rSkpFC7IGV/9hME1Cxz0qHIzhtob/rvh
he2il+DshH6lWSwpapI9TShCuecSyI2Zc8nT8buN7LorpBPzPgCWRk0U969yNBOa
RsDLn2zKRtIGnJjWeNLU5Sk+55UKgNHoDAeAXOZPmOgVegYYT/YIEjjH7YQIwB8E
4lJOKp0j0JHs2mTBJe0kpmGhichHKT033tFu6YjlbyOUb8Oywv/xEbU0b3KfrXtZ
a6Rwnvg2aD/O3JyZg5W12kuXqhWa7a5w/p4TFbRvCkHhuNfBZ7z9ZcLp6xIaWw6i
kUzLXwfNZAfFiqJLfjFzQAGT2DHqOBHehscGRZtM7mMtSUjvnl2aFJhj9ZreO1zW
6DviS5BbMXkB1OYpy2GL6yBCUTU4Us1vonwzDAmZgudb4ROPNxfbCrG0hkmZoKL1
nGAMlqvU5gbcRVUmwAO78+8qmHITJkdY8f1UDggKYIOqwp6MsPMVrD+9aV8XYU5D
yiNSsEO70T+GoKO4Ex/k8e/FV9IHXKQjj2mV7NS25+p0B7x/bfG01PGN1ngtD8Uc
3QqebqOSvt/5LB0DzJSZQHklpXmHYdQVobzzlQrQxGbuoP+AIwAiwlVq6fCNqord
28YBhha7w9V6w+37w7krH2bp++p7FuuOIZDjCyJzfQ3VwWuolrSkY9iiPUyXavzn
JVGEw/R7kBExoTj+pKCFetE43LwLZIonSf/CiW6XZeGoonjFwxegOZinkoWevGoz
DqR/5oJ12yzsyvAiwsLhCAJt1W/ibcUvxPnFyJUvXwz34X7cMJgTL9ynSlx4DQzO
s+Wrbq6bKA4GagcwAxk0G3HwLhv2vBYIK4ObYF27F0Nfii+hIrFzEMQzal1je00C
FKMSXes4kaM319ISUz/E82v2DurH8dyl9cLCovDz1lCBqTCx1MeOqD7iw3ZNzjLu
+3LxsCS/0kEx1EXnqGHyIiwsHalLyO8yVDVcj4f2LYlfEyCkhpe2m0YfxUUQSVz7
S6qQB0Yp/CU4fwTPLIFXwO0+rqtAOWbpeYhFmtbiPTSPMQ5iYP0gg8o2PmrRaYTv
gF9idP/OkDjkYWiwST1Vxwk2TqqIbrmdWhYt+42UGHP9aGVwJ9cSp8TFgpzh2rRt
pMvYwXIej7SgRE570s9xI70s5M7bw+5hjlnQY+zp1PE5l0jndu5DarDexSeIip1B
usqAOssVIip8zOXlK7Ov6aQgUoyiTBbn+zmdq+Ygj21lv3z0lo8tFT6VX3XaT+mL
IkRXPDSo3fy7vFMrLlIrIW/0EyQCaXDFkF7kahSGGcXhxNLI5xTuqf/zq6m6avyT
rFRylsZzyWinYqmNcZmPZjeP3jY6kfYJv7XUBYeFdRletycImow4qlwsXAMmg6aP
+HT30eKYZH7Tux7ebNRMHxEGn4x4D+GJqjlgpVHRSZEi5AchdOLsDZYvpZPFFAY5
7EhQA+Lc4SO+Mi2TSDFrH6s5SS1xdeFcAeBqbt7Q7ZYaAcuSoRv7Jplg1hcaRWY8
nmoUK50T0Wjqk5mQ5nTDUNXRGYNPpS0Rovj44gkSeJtUDNqmSIFbyUyP7hdkCois
TLodP5G2V4qyqTcF6nGXDzeIjvrrGJ4wt0yA6gjfrHVmwEJJE//++UW4ixYcvGca
Cb0jUct9sDJFFJ441VF6uE97SH3WOAUgx6iJF1XaPnSIUO8jUiyGnaN7Ync2sWrv
y/QQY6SqP6OGKvXIIpYpe11KAhgXjiHcKHwlGmtsMG+Piko2TAq5qtFVc6TMoY/d
J5QAhavtwG9BhauHhY3WIcmQwTPgikdLUjTuU1HrWuArfZtd1YuAaoFZVTOX1pYx
oJnKhCC47yHD0uwsVaA7N7tR40GJtRLwBawDOFVMrispNXXoQcPCHeV6jxsj6wqs
ORQQ+dA1S3hZ92yzvfopshFGn/AeuTEKi/pTp3Hdp7SxvO9o/2WxY+D/wsjjq005
YnA75p1kUmIgLQ82MWI2osojURARhNlbKv01VHf0vktnrlKZqwIKWwIb/fH2vqX/
Y8SfN9evfb0Q3sT1ICYUe5ABNvrmt6lnGJWnV7egk+KXdL9hXtUoPG2i3lOWag8c
Kh2hz1Nw1M3PwQJVyof260KHAKBrAVcL3sgLXzUu7fAiMoVnmaVYvNk1vM9VIiyb
k1ACetUTW+G/3dkb2BOD8T5orHka4aMovTtHq23uqr9qZHTIJhBDuntYSgmIVflO
uVi/4OWoAe3K1EagXpdtl1NdIXKTmun7dRoXGJoTDVyFFzO8hOGbZEWsP8mMnQMV
QnPr3EJffA4DbsVlk89xsaIrYwvcgb3msbnIAewvH67MMnGc5uSsR99M0CJ0ApD9
YG4OcILgLeRNVX8iMfLmhYakFXQU7U8zKAhZkpDKE/OHObEPRDOKoEJsmIot8nXT
lu61yHDOgn1diCvHPpRvuDimKLoR0rwda0KoZL5znG5g9sLJXP7rj/G8JUmediqw
PU9Q/O3qIVMoEp+LBdU1jkQVT+ccO1Al5jSoePmNWtQZ2iyW2Ml+Ao7OLmdDxaW5
ZSfmv/yawmjzs09N9JzfDCQZEUC6TdMLLJTUbUYeodzi4wTIpmpYVOXdab2L2E15
2VdVV9iZAFeaHq8HNMnipx42BCqAdFG5jEzcKEtd14BisEIpcz6SJdMaFKaYqRGj
qXt/2rnSoyZfOM9+Hu+IUgBS2zvOA8sFzrlZtezq6MskEQXDHcufAOqRdj6vGxOG
H2Trsdgaxre412sdxJg1qMOAuAmEcGM2WcBJ4nn6h1OxFPa8jDxEE55zDHKzkGj1
+XwQRThtFiptCwYljapGMKOf2Rpe869goY7D5DD/R7Px/geJXQfDUSaV8ID/eu39
DnPxfWzHpalaGFDSfOiBTmqS7njfPmxH5iuo00nN7pGIxbtXlx9e/jz1R7XVv4/c
iO+ty24zLaDEfZhTneik57cmg78WbQJaeur2TEUUSVKB5Brf1jk+CIuY9GPDtsU3
zlMB6xd3RbjAekBxW45hijscPVFrRqbM/JiS9qrUlYPdTFbHrw3AGqUI033OUfWA
dxm1N+oVuUCFm9S5eyW/Bb5lDi1x/GeNN7mp+KE+DFkUjwNafOL2vMiHhC1a4p2K
uB8XPecOkzymdhWqyg2ELSefGfRgHZiLOgncpaKIJajqo6PHIN3MtrzXIFY08olc
ULWHaOeTuQUcF8oY8askzVxu128S4ChA0S9L/s8EoPrNFUcBlZMwQUrWp8Q+wG+1
b12DQ3ipJRG3URE4A75PNtKvbnR3ucca9j5MGUN/ZDUmNeTjL+7KUq61wDLVGpYK
b+X1RAK7M04FzHHtcZtk5Y613dzBUdpUmTaLrr6aRkVwuOarW8Yqo5/pPu4PVBOM
+G3JnQrVtImoS3ENCODA0/8S+RR+5esf99RVuFMBfglS/5EwHsjexv6NKS1RFuYF
y2Gu/vrGYpdm0POjZbdaZcogbqW3KJH4SS1037V6f5QQcx1FjC6qC0qsVdf62Csw
U2CJvNfwl+2fCnKkEiwwsh/HGE3ZOUuYgjcc8WiF87Qz4qfwy2nXrdevA6EqSo4m
PoemnZFljYvFOwvHpHoGXbjvXKBSW6SGUUF7Z/ppJucXriLSyCKJ4/NauMA6zkNG
LUsgDiKd1krDgBWmfaYnEjyIpUhmTbYsn6Wo6Qgvy1vvZlcRseOf0av4U8FVzthz
QwY9YfJwxidk7YilK8VB924+QAEK1xlzpIsXNqhVP9f3BK6XVCjmgPGuMzY+Mqg3
Rd2yUqLOrFn7IJAePDHlKFi4Qvr5RzjiRqWP1QULlsTzvDXyy5bWtsQQRgpDKBNh
hIfVKUOywuJo7xOHV8BbyQsdazYRxvRvcwxH7SzUe9/sfT8AglEW7Nj/rjIKHa4p
IN1tGOHUa707o3cf2RlXJ2MJU1lJlkSpY2LJJ9nYRVx67VPmUXBZDruJQ8swSPtq
dhlpDIskseWWefzYDpoI5esX7R0jBB62/rW/IGKHZfZaNS06k8o3wq6KRY83Rtbe
Av4AiZtD39XHoom/l5ztywkdcSlHs0jQDtbgd7K8EI0J33+SOHIHwYJ7ktnjv4/0
MSuGFb0my6uax4sjHdMK4AfFi61PFZo2YATFOaTD6vTLxdJ+aVLa+Tc39XioHdwB
KmyXLjpAm0AKmItpxsiemEEOxXGlxZ5w3Zl8RhEXQ+KEuJwbIayAmOgoPZPWHYIe
ngOfUOJ02Hx6UefR/vGL86iz5hM5u0T5gacypfGhWj3THzUXkXUvj3ozTzYm2f5J
2k8kMj2eWTSWV4ZHjLgDv96HA55Ac9S+5eDiQFtIbP4rfy8ySvqzUqa5syHYUeq6
nJgfBQAutbII0TitoW5LWdymnno1IHx3oTAUN4uYViZIo5kKWSyQNC0FKO+4xjCL
djs78rcU9o9AHD4Embqea1E+MNx+9vI209gOKg6H/k5wK/xY8vw5GwvaZ9s7h4ik
z5twwpLSMB93VLAZuLUJCK5i2V+nY7V79JZ9CsOlelV+xqDDjpgu7LRl5Q6fR7lX
fAU6rZa0kZEFjR7yGIa2vrLCKm1OMpcl303tcT/wZS3JDt6U79QsxGA7jXscrrk0
nJHEXko9QZeEBZDCjLUwEuYt/ggbMSIevhmdN1CGGgm0IMaYypw4t7c2PBm4/pPi
Iva4szpsTtCUr2Ocztdmhy+/+55ZFBMTovOAVD0ZUP0W93PIUkiX8nJFxgv61s7b
Af9ueQk7MVZ9H0vDyJxZm8MzMDELfFfjBAw4VqStK+ltIguCW+D02qn4dTpgKMRy
DMvWGgC5sGOkq3hboWc8iIS8RorOmwa8pcYgg9BlThMaBZ3tZVkPwfmnOYx2wtuP
LD8gdKphUobhSR96Ys2U8EkRm/B8KJUbKOEM/zH5/weaMCeC1g4Zgy3eUWWH06Ql
GruAQ2c7qYGYPP8NQqfxtVXfxylJuhD2aU5L02ZS0T2bkpsFohTQLqtL9I18oZiq
tYgACYZF4JE18dzOX2Au0geEJZ9HJBhenOqKHFRBgPYUS1JQ4pMBcAk160cEDFDf
++GnYpXA0lmu0KCZmMxPAur3IBOleGS9+6fOA27mHRqc0id7Xh5drKlecuowvQsq
rT8/9tnBchnayAK6m2ew4wqG9bp07x3ChcI28N16zPJaIX19vzdc5DOjNnLitEzD
p2HKOC+btVjQj0QJ44zaVGvUM9hE3XALhcNIEEXXYKJSk9gcn35rqpfwcOie0Vl3
Q3CNusea4bQ5oDvJNYNH9pFEi7+H4F8VQSYr69FtV/DL7l3mlDrVVyWc+R5qLbBC
CDiCuyr0blhsPz4WPhUM5cSi4XwDCkcUydWtZAXWHJdc+JbJOKWfxpMioOMqhyXM
267vbeyQwIVZTy23aBhkvt/MCC9FkBCyFi94Ms4oNqSzA3tx29ae5V+bDvU2JuNJ
fN09s4OdNjXxzflacLf+6cPProRr+Yap7z+Tx8afo2jB0RvyajeZthBFPw4nHadN
zzhzOgHTgLG74qV7fQpCVRXzlKu/CzhFx+yEFL8kTTfv6TOqQEHy7YEMWowaLo+T
ZFkPuaXY0oUOPSAEFkyeeDJVgrko+LJhktSnDEFUu0wtxY0veCuj4/+lPtlj/zN4
DVhFxqBP/l5QvcN83KmuWS/MZfyzwvs7gsybzzm/XRdhUF2qS9B5lWgWUut3MwJq
oRpMjw+brCuwDbf3CIX7W1xbWeEfObQNMqH2dQT/k685L2RIceiLR4gTSyr6H/1R
MraAcN5h+k7tFNp0gRgu4PrqM6bY7OJ7dtHKL2DlVvaDtGQMPJZb91reAz4KOGOZ
hLFg8yClIge9b1EAlLkF7lgvMnBhgolbCWvuEsd/q0wyf5+o14le7j3Ax2q58eNf
0oJzncCxVijMufmZp2Mf7K4e34g+GHN+YydfNYbedsD5Gi5GlhRUzBPvAN5OKt47
A9rGQ6B8p31A85OBZbkyJWoyIvzPTp3asc6LtrsOm5HFh/2A1uq6nGREXC1NQgev
ZUV5cqXVqFRBsXnQKwNZVTAkKvHNIw/rcrQKxO49NPxIEEav2FysH39SfPLeWxhj
Aw1bIfd2461Yxg5Mbo/kKsK6uKb87MPFHzKY/ZdF8nQ6IWmredCPz1wjFnWGfx1d
PS5tZoX95imADVM9Ey21iMp5XnvVu0/tBH9mks4u/x5hYJzKh9xMkogVaE+iZ6lm
4poeypn54rgyo+wvriPCSUvO/FEH08gKDZP78TG5iSrUkrjAkzb0J69T9lRmQzZj
p7g796l5Oxkh+B6Z2ycZ8G+52+0eKMR1B5EGSsR1hsTbx8JnA3+Nf2uJih++YyvM
KVvc46TwNpvMCfHz+amUBbEokorQ33Arv1T8+7XxDAmmdMisyFAqBzaNUj+S7eg4
Hno+yCDfoUyRZ/bX2MThE4bdEPlC81Sm9+qJ/RD/sUBRWhBvhL16lOzNZV5b9D9D
6wwEH69MoAyiC1EsSWY0WPau+xiEKfD5lrlUKnKLckE4L1XmBGbK+1p+vGFcNkCE
3mCT3QWdq0oRIKCqzNDPF5aXgrb4TxkMOOFami/wjFxQKlwRSMuOZB+HdLUgrQYU
s4CRN+npSsoIx6ph88hmMJNWPGORLe6FlQGhOEpQOYhZtThetAFqYfj8X4THiE9C
TVfo9XQRKc+yna/nLL1foFpN9+OL40gimJB6QYpvylRhVtQr0uj0UIDLxfbcG9Td
XiG3R3+02fWItnjpa7bXm0utgbF+pgiugAqR2giV6oClT0Z5otwCGADcMq7BMdxO
daEMp68TednrGW3Rsgq2QmuSLAft0Po6usQ+fP7vGlcIgO48JhPT8b9MKV+rAJWy
u5wdkCP+E7KeyKL6Cn90KzL2uFHUHXdSJC90DVLnwZ7A1+hNKt1fWobm576SYd4s
+/pDNsqj/IC4xrg0JdIhO84PRjaE3loEGWC8MWERC6iZiPmfYsoXtzd/kQQly0kG
GxUHD+0DMeqkU/4zgyj0NDyNjx72P9DKTfFk+wYy+pTPJKiWPawBlk5rG/289xtY
w2lSaPQRVdo6bZqAzZ3F2obm2QrR8L9TbKkiUxMwGbqYmZ7lTAvZNWqDRUaxcqIq
G+dq10oiclWBOgC9sZg9LNpdo3bqb4o9/a9ZP/FyUizaCDcgoJdeZ+e4N369EeUa
q11pqch+HMACDv4pInHv+0Fxa71CXc1gu72O5pI870Ubjhb7dU/7AGIQUXp926HF
RTWjXBPt45CTkMJGBKBQtZ4t9aAW3cuUfcswc5QJyXXz23Na0mUTmeel3GX6R0KX
IoCUEuYZly6ImnKKtNoKWV+H5a8WcosiBSnl7Ez6LaZEwFm/AeYEc80JhA5ZdZmF
PoTV+/UX6KJf9NWFiIdxMEeulAgXw0ilEZOLoXX3hZJAc4vQCb1MZPHdhuXIssJ/
7YvjN8cNa3i5mAZ3TgQc6QYfJj0+H7IzC9WW/KB1rDBY4Dvnhbtm395fGuYRa3KM
JHyzm1wIENQL/kFLmU0GB5N7LzUopfret69Z35N0/Rb1RAFougX7Z/CdvJjV8ChM
yGHNr0eG+/cQVniJIMAN4IluvtIYIvYqQBcXA6Za7nKctM8nbjTasz9qxI2NUTVv
RO5sU+jH/n5itKYkVhKhJjHJc0kBPVRwqgKJ5+VWgkUyHxUqwpiZ8s2v52hMeHzy
DiaAw7a4VQgv7ncSm5syxSSFfAPXaoFziwLAA4yOXC2qALcc2eXUwoKslq/3v5yh
7/3IlQODBAJx9UKmJUB+SW+NBumoxtM620+w59uCJkFIS4VXROmmkQcQGpc2ublx
R0/KSu2L4J3Wzf0oAPGaDNp7QVNCP0HypXPTo6zb4vNQvVK8d1SCd8oQXakffbNa
MWZglifNBC3GkE8+ib38bUBMfSITOfpGfzWSg1bNldwaxt7HgVKwZN0xWxWRHQwZ
doeeJcfiAL2NLWmFkL6ZF10BFCB4EnmIp+DnbOVa2wmEQqOIR6ABr5qfhrGNNr+z
qhNORd45fjeQmyeAZP+IIPb3JLVfiOX5IDvfdfruj7HuFJAd41lQY+U9sRekmSyp
N36PHiJcBu5fUdinOl8yRKkBOPnuucS1ZqWEyRjzx8dSqZT92ztA4soO9MtKudws
C9KAhoH1Hhao/psk37wwX0njMFLVQyRoWRP0vBh8SXBc4N2jDP7hgESPHLwTqpjl
MdklUZPpt8K+n4SsegXYLGkqjwIdWGaL0bIOPsYOdIEXqyK7tL1svyjcUhukM7YR
2ibySNNpzCikE6JWB5AgSuPngbWvrLp2tQMcuUmUTxbe4IPc8xJlPlUSg7swpStA
PSxW7lGqGailqIiYYVXYwR9kXPSixFNxIb3B1p83FGqYilsPxeP3KLhW21AcnvnK
zrLubCd316kMbxnIhit64oKUdSnvlWg4FL2c27ZZUr1HAOINto8DH8/kiwm31twc
+VD9lcmip49S0WI6MnH2S6JPjHNsKDEnO/k1EDXjepTdqXfUGKzbilAOUFjOH9Ty
lO60tk8rxME3jWmhMNbqN0oVU6venW75v841G46xw4jTjmB/l97s/R6fw9nkfpWf
yI1cBxHryvFKVeAzekQEchlIF21USzq6nKwfIqoA85IcKtgUXNJY9KwiXpVGZqD1
BDIdjguH7tLDAbChSnW10VUjvdaFfdg5MoefQCwnA+KEUNh4QW/AZFxAXWMtOBvd
vQlW7u0FZ0V9WxA5cMxZADwQGir1qDsWX5PRZM7/0m2l+ftZATve8cznYAoOyMos
WcyvTGzGBWt0G10BjzvgTZvxfYchHvprLaKTaq14SF9PbD0gpPlhPEM3FsnUA1mf
wmW9JbQCakMaHa6AymbeTM63YBuIzZnQ1UUKEWtM0NxU0TaJi/cMkhpmt15e8A8c
inO74De4b2za8psR7PLx6A==
`protect END_PROTECTED
