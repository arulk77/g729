`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
D8T85PipH0DsbWL9TFzsvFF3EnPRcj3MvEp/L1+X+1nsXR0ephPdZBKFtG1CfLz7
3p7VBrke/3MklIsODN4RDosOirkdY7vEsUc+TtTaBzxK5tzJCclkmzYExJzayb0X
Cj0z6nP5iBKddu0e4KvsIHz4rmloKwzzZvJnQBoYvrRAu6995QarzeWHt362WSHx
Ysb8LHPpw36dMmzst8W2q/Qr4S1iuNDsVj5STParMB5bZFn99ogy90CULGNFB19/
DgxM2RDYBaMWyMw7fHiGqRQENjQn3aVdUWoBYUtgyufGKZvJSP8aLphlImFcN299
raN2wYtU2l1TSM49MYUqJwwDhX9PtD07PhrG1PRMn8dVfAHMOqj8cLKYplJKo4mW
NPghDbJb0+NkH+8R8LOolIS03kvuC6JW/lFiSzPNsEomPb3glaNMw9sILz+bpqFd
YXsKSgZh/XdxCgpmYLr6uBAT5doX5qSVc/D5HG5LWB9fwJN6XzU0e+WQoI+9R8RD
hVex9uGzWP9TmOlMxtzZGbfHNvXToL62WUnMT692zih4LE2OT2jPotMmGG/Ksp5P
zGvVYMBfNjtzqXzs6YhaKGfyEYXg9DuLtp+5OWV5jiloQpimzHS8PFHO3ahruq9P
fX1KpqsbJDZjDofT9Hwr6N7YSKVSyuBNIHIm6kCrStZgKrpVQobukslwC1oNLdEL
27S/XOs2fXiUXRd9w+6Y8AHcsxuHXN/yEqatfnzUjOhPy3wPTrA0K1PgzD8CIH5t
yVFoGa53rnoqGARmERWTvOQNj//zcgPBG3Fgpfg9xlPBnhCezYFPoZ1mgllmCHjK
/a6VJgkNX6sHxHIBKwwVYrpAzUgswDyS1jl21+vuNHeIppyNIGVP3nh/EhXHt+D/
jVSfUeYEv/kScOzjD5+SSz/qQg8R/pcAZ0FELR8YsulrRGqMnwbUldhpMnOzL3bn
1M/xk2huZ10NIglUcqDUuCdABze/xssEGIGEkjizew3eYKgnVVTD3zDqmDcKWO6b
dERM4yTxz98SopDB1C9DDIZkoud3Bp1WgjS5Bs5YcnO3+/Xgq0vwcqy/DWkQ+TmS
YBkQpDBUvQsdgBMhfGlC0ouQ8ACHg4mOlS2uIyPScaxByi0R6eUK4rCRTQrdIV5k
52hDgsoO22JT+Jka6AAsLwXrqu4NCcEFFXWXwAwk91djgG9HOdm3XvJf2jByzxHl
4b6beAaFK3i95sBwj06cHeAbNXepGIcRv7gXon0/Pdu7cUpr1U/Xm1zcnHKe1EyV
cKTavFbYNnU9U05WIH06pZquKbxI4YVk85kNRCkar81N7IblpcNdr8m4mFZHCClx
D+i8QaGWFarO7EaDLZI3LR6bJDoNaX3AxRXLhzoqTrz7cE9eatrp70Pw8x2Hv/eK
WHwKXitk9CvqZyt/jDO/nSYqjXc5Y73hEcGKIOWPkn6HwK++MyFf+QTJdzieM5wc
VFIVVs+Re42C6szAgoV2yEcLo7o5Z/ChgOjWPbij5UxiMxdvU8ElzjUaSul2/un7
tODGU+CkAHq+SYSqIvLo/wbIqhgi8+89k5jtUzNbj94FQWqcaXaDuVjs23Y24/y2
9LQ3YnKmuaOxSEBRc/B0UAnzrGA96G2JNWykHHkf854leax5MQ4ngAihmiC4502J
JhdRKXdOABWCES8xA7AfjB93ioklpL8f06xkfo9saU2ElekHUqOryVWnfSnglxIp
qipeoY+u/o6fj3PIrp5xFEdcTk6eFNIgsZilvfV0/UFXJeKh9tMAtA1qzjiQ9+Kt
3ExwYB4qUvuA1vW+F1+U8T3IRQBfJVh7rTr+9YaxynXNPFpOGvyofxW2I3M5Sswr
orlp+aBj7gh4cg1L5RP7QCrrjbttZHBvtxikxZInXefM9XNzs8MoJQN8NYeSQNNC
jc9VeVgx198U7qY0yck+P8AHRk8/qtEZK7FzOvOf2hJg771JVj/CktUPueqKG2aV
zSIgF6BmnKMGPNzKQT+EEo/pIufQ2+CBFkG8RLk2oaIkoO+r6jV9mQrN6Uzx/b/R
Z3lZXhdbKY3/Rtyn1/yF/tm3w+T6ZenmGM9KJHhJQvvceGANrbqaG2bSU3v1F2hd
cV5MbkdWUtSi6l+SHQzBdFkDYYxo2xuDqJdqf5Zg8z4CkMfdJPOaSsemO+mGbTRU
+Y0mOPZ4Jm9SHdvjK5aGWANjmDCYYvYJFg+qV2mXYYQpbl65inCPe0hojrA1txBF
UuU4UeO1JY6EK1VtDLnCTO6eFrGAB7eKWHQhwHBByJHek37fKvmqzL56JH4rmiVU
NhB9zgsKBSrfx4cWn9I1EnoeFBWB/wVuMHKk4kdBSge84YjfDzH1umX29wEdhl62
n45IlAVPyXKGKW+u+p/B9PQSs5Ph4gUEYjVXCdMUJNh2nW7pHSVCgwGrkfcV78Rh
O9utNGrQLcMxqrL6TOaxuGk2/VCxzzObDrKjlUhYShxQIVvdpch6sp5RGGt8snZK
pFc0ylL/uN7fjbzPE+R5WnGzNdXLIP4oTur1q/QJXzcJimTJTP3pust3mxGEx7sH
damhN2Fer8L9FC//IZR7a8rfX0oR7Usm1kPE9lTvTuKdpqgZy8ffVCOneyj/FipK
ZfWBJCY0k4BUFF3f+3tUnUQwZSKOW2rA36iPP7kMOUAuQ6iuV5Vie2Gy47vFuwn7
EvQ/ZmSwYrwET5JZS2e5i+/dDeYdWz0eplwfHcXpdFs564qxUEXHpO3w+pLAGFfg
hfdU6j2Ojg2EhXqQAWQWVLsSqfdAoVMX1vjvGvjb/A8dkieXGQwM4yTtnFjL55Hd
JVXuhKIFeFKBabNKLpyo7R83u2Cm956yQUBR7EcHFTMUVgjaeuUHJ+2Bss0NFh6y
Awvm8yNewK9PMS3gVXwHEjcd1zdVqnKhsEKCUXzVHIm4vkPypMb3ulBYXVg12X+1
giJQq0m3SIVtJuJ5loweO4BhO8i7OnVtw1eGoSV3IVjSsWruKZHPCcrGqifTJ7aS
19k4vb969aD9HTzDULLbIINtuWVaK3Xv1Sryi1TgHal1HDdbn//rh5AIBkDVFPMj
KqPLsGP1b8wd3uW3z7JLx/MpZZ3JEXVzjIP917Oz6nU2/HJTi4TR0zYX2oSLO4y6
wnOm1dcROTxRK7IlHNlqCarrbQ9Y/jPgI0fvBZenJ9H7js5EHD80B3PbhpZnLfPo
jLg52xQwfyYmF/faccaH5ouy0HVyeVQy+KUhYhKRUHw1Qm5fUzBMaegEs1hTX0QR
IuHD90OS7ydCt75mRVB8SMlkwmoY5Yyb/teJ0O4wNKN7KZqoV20e2Jof4lJAvqrr
gg3qyWI/pEXxfLa/d7TUtAileN0n4eCKahr7rNcH2z0vvlVO2Q2VGomskpvUC7B7
iy35R+qShwKf7ZDjt2DJq1Bq773QTZZzN/n9xTRKURDUcHirYqWXaX4EfEq2kooz
gVVlYmVoOIDljb+8afcZr7C6vm0QQMOV4OETbOT07bBNRy6QvTwSniTS8WYx0He3
t3IpcHJnw/ht4RFYm1wj/+k1BDU9WVhrr6Bnt7s9pTyy6FV2p94NFTG4Lxsfg+RX
PtIwiTHKxyZ1p8NbpOyH/UxvklSR8IlLvVi/95gAQQEmMxgxGcPRE/EljttJFwam
pm3vNq0DxN4ptwXiYPa1VypohZu31F8eyGa4mtCoNg5o+i2+8Kqg6O7gs+HU1wre
`protect END_PROTECTED
