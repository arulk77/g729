`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46s2eIKYkD/SU2UBtLctagWd7xornVfkM/rtshyVpbA5
oeol3GR3t2gLakt+e1aVTTK1xsW57wEcUI1BBHjWyeEpE/vBvcDMIX2gfRtkWN1z
124IKXTrf3eI3CsTL/sIHMytSSbEBagLFIXITkIwFLWKayfHLWmHsZWqTNvsMCek
BCzoFPqamHAiNVxa0pTh1YFxNIz2J/2OnKHs1G7ydGS5Dzps24y306rt/zcMKuiP
b3ZZXQKN0LeXE9fqP6Ouvyiu4ejMteFElO9zKWzCyYnqU57WpEHlJAWpnl9IX1S3
vfnV0KBcyDgwOpgJ8O757EeBqVosZ4UPh/EklWBuaFiTmt3gDSvPDdvAO+0H5lQA
FGQqsjkPqbcXKwxXeAe1Yg==
`protect END_PROTECTED
