`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJY7XJiNmZokp29pRWC4Wo+GyLjMatw+Srrbu41/Razr
t2+Fj8IPXq1Vq4io7/MuJqaDdSc5eVjz/T9WPiblIoZ705LFE0xGfhPnt45MIbcx
h2IhWId5xghbhPSE8DQN4IQAWqjSw1xw/GUr/y3czdblvRHaDfWIUAsVtXiFeJtw
pmBJJ51v5KG1TOryZQPYKpP/0OiIEqaatzc5fiwccBvDcX3wAcregplfJd6s1tVd
IlS7ODcJC2MsiwhVQa8bMcMhRGPXaTEbe3TZqasc4fsYwzhooZU9slbLUPzJk33U
uUIzhLn1c4rlKPWxOI1XQGsmTRBDH9tnrMZBgzc0fOGGW0Fiw6mjfmlVkktNxK8N
EtMUbqYt9LDa0ZNuNTfzn/m5BmUThnUnOZSyPw5lXrPpJ8SMQEKDUhsEr/HIorbf
k5dJ5MY6ajY1+DRM4L459Q==
`protect END_PROTECTED
