`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lu0QNEIQtX9harzTXcf5/YgGUHjI1qv9N2ffd7xJ0rWTRRAM1oxqXasSNa9uPfLj
JxwBJtGL/XhXBZIpHanyWs6Y8VEZmxo1uD0FXI1cvzwA7vzAUsZNbVEkkP7cj0Su
5Z8i+4QluRyuPtf540hp8MdSn4mnvZxqRjyNtNzSW0gbU3NXW3iyRpaGK+QqdFlk
Wh14Am+dWQBRcfwXI5ww6pwKCmRI+8heCdIUa5oYAlxeTeYEF14AABQMtIVsp041
iIBi9ZR13uu3d4L0DMHzgaSdEiCuqWvqfZ24O9uraGU=
`protect END_PROTECTED
