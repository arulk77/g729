`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBbvf13VRBkzEnDemkTrxKwjwR7rPQ9DDx6inA0nU4xx
Osn+9Uxq9qvk8ibRx1kBPsqucVdXHAN+xu2QZI1VcNqvRxRkbuK8pWpCzXFdu+Si
iVYpGOjM6jYx72jcteevQDpWoBYXcot5UPmIUNR8cZX5AsXTQHzt0gZdLELwNqMG
QU+TCmnk7qGnEBTZYb5xWSF78bas3r6Z9U01JrioOHFvzyrjozPN4VRATKpOk733
`protect END_PROTECTED
