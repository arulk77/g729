`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCBrhFMgiYhRFKq93gJpyDD5HHT8g3QzDPY8WeAshHDY
2v3jz0QVymGhKj7bIAp7lhwQozvbjvlqhjliFqjVfGgLrgN0q51+1AIMQWgy4hB7
UGoLAWq0yqFerijIrwTk4D7wcUHXWWsSgoqyUkgqlfl48hdotA+TR1fCsXHx25dy
PP3f/CpUKy4iDIF5lPYlT6n5waabVlQGVlTFKziQToQmqobcVarQkLX16gXNdbyb
KIfauNJNW1sSuLQy08DqaUXwflsz+7uAj1HKnC3wOFs3PxdKrJTqtt+k+CBhI31a
YOa0Kh+1VFzG9vySQk9u1/21bUdstcL/oar5YrqXHzNIico9TQIb6rlesuq82i1T
jo8l/010jmFozGmYjBHzSQwA6dwBfuGtqpKu4GXs4ZXR6xu50xuud/0TQ1iA/yxJ
JJpb2q03X4WeV26J50ktA1EKS/4/qlvShM/3HKP1qaarKSDXvQtQfvYbgh4F9fe3
`protect END_PROTECTED
