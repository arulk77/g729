`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Dn52KkuUcMNqr3e66pwaUBaC2CYeJsfRzXfHC9OsDbeDTK18q92Xwmc8yoNsvGs7
Y5GOQ+JSMzjUZS+GoCFvK3HQ76P8txDX2M0nYqnVaidJOiq27MHSpks9fY3rhTWU
/Mw1IFV/COK8zG1kQAAAXJcHb0uln5RtKQWtNe5RMwuKfRbZcTX2Wz6sAjyEpvRy
C1EdcrEOKug3h/ngUuV6mLcpIbk9zCFFuk2/g5awYdbkdA3/VgrDnuVBzQgp0D3k
`protect END_PROTECTED
