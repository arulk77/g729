`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEni83p4PUxF+TgfY57PxMjQ9ZO754JbjKripJ10oOrx
uv0QlK6LKW+sBxHkAC6wr5K/daDzx8a1j/TTp8Yl8XzltbxYTxoojlrdTWEMJUI7
gt0FXwvkEnNG4MiIF2jkTS9PgcI1nV9Xwm5neJHCGO4Bq/r9YQiQb577FY3pFKxj
Tg6kVX9EUeKYgx5cCXzUGd2SRTKkCw/auVB2jB0vkER58znO2WxIrRZn/pTkX7N8
22qsK9MrL2RKe3C8AeOPCQ==
`protect END_PROTECTED
