`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+j/LRsCNjWLGrKq/VrbLK5kh7pOk/+D5520s09jMFhZsl
xiG1iuGx0MTndqEwtUduPs1Lk+hCkQkfuxRm5IOLtUj+u7bqtqCBySmA0estG+84
NxfR+cVCNp6pSozdaXt73d+8h0eIw6xfS81Gbuja74VVb6L0gnhbCA//wtPybcCA
`protect END_PROTECTED
