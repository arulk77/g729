`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM8FFkBYcpgabFKsg0RwYsLaJIgNT8YSikrcSbSCDutV
7H5bWKdamuG7OFnqes1pG3ehrTDd9MZIfz+bkfkXkZiZTxCbqxvlMoaxftMjUrRK
Tyawl545IhCzNqbZr+lfgueF5XLOVQrWWCWr+fCmz+SgD6e0Bsc8JQRdGespRlLe
Po8TIolIba2KQQk9/V+epKii9Odq0e3zuqsu+BvuhGNu+K7/qH2ORMCBzkb+3Cky
`protect END_PROTECTED
