`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xhzHJS7LiCuY4ToMPKYAhvM3Yofwml695yVDRC/L5F7
FK/3sBPrcrWgRpHxG3XcUbejQ//VtZRAlsnyoCJ0Tkp/1+o9K01e23kWbLJF8KfZ
1ZCmiyYrzKymrQZf14wQrwvT95Ynqll1LH97GLFCSwUOIglBS5iZQBgvVu5d8Q27
xsX+YWHvNRBYJbSLvAVR/ze96iACx1hTuqc0R4I7WYK6YnrRQ4KqmnZSZBWR6j8I
4a36TldH4YNLmbakxmqZNOk/WoJFSbiB0K3Ju417DA3YcqtUHPzSAkh8oJYnRD0l
bT0OyL5mXcXEEqDW3yvY3XfkXqruXE6G6wiDacr/tDCTLA6/nChcS41/EiwICMlp
Kld3xRykA0ttBCVq+acmjQ==
`protect END_PROTECTED
