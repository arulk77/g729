`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGq0NVotRSGhQUx4Z3c7lGdljl14e8ccv/jzqlFJAzgP
WKmvCuWEmjl108UaPNSDW8Wd8KNDMff9aXZTf2269YMAWkR/4ZPNclxwWOMJarX/
U1Va+sCsV4AVKryAeudgTdJAdVgVPP/zij3H39T5TQYN9WdT9pnZMt25ilnIv8NN
VOAh121G/PG9WfF633KljUigXZlVBE2wWv20vqa/wNJlSSaFj4qw1nufxaiieiNZ
NQVbzEdLrLKT+txHfNKTbhU/6H/+1uCwHBxcx9ud5AU0B21jyI6UmW7qtQO6JYaT
hpudnW1rTZDaGnfGk6l2wr4czbhHktZw47CHxQ7X0uFJenwQrlPvG0+W9jPEX+Fv
f0s8X0sE7h/wdzwI9nFo/vZ4QTiseImRC7xYsks2m6J4jhza31EgFOm8K4YlsfA1
4+vCV1WO+5nUV5eGRjJwYLdcC2ZzKptz38QM5QGiqnCpltCwQZSk7f3E9Wn32KuZ
Jxbe5t6mMF+GN28R7LONy5Y8f0wnHFdvF4kSWiY9HzVn4yrhMpy17+DuovqX1lqN
`protect END_PROTECTED
