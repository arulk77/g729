`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOz10Q2URn5x5LgK6T3cabDVVuC2xUdHkaDh2WOzHWjp
HE0oMtmuW87nsV4Khe6KAdwd1t9QTlShRjLzBSpG53FW9AykBR19SW7z3bwerDQU
PbqSQ5MJ2geluXE6xHMO8ZCps5vJS0/RwqmhkrXWWdA8RHUWcCdqsWGi32fE2/EA
zCKLUgMS2qAH4SYP2+Ruh5Ho+XCUAHbKD7f5SlWow8EI1V1A6toNvyR7dd5xu9+/
XGqxMHJScFGTJ0TqCdRPvg3xnHiEy+kt81fBZljwVXVU4y9mW/6ctow9FpUGnCNm
tnOU9OhU7LcPC7NRO8DBLRfW7jC+taNauXLOXsLMIWi/91DRjA0KgZ4nwLH8usB7
e3TAeBaQMpqFtqOMsojWE/6rUNRVA3JuiXKOIW2uwmMIkhogF08zjjpnMwC7n3dg
BibNMC6MTWyjabQ9NdxCMbIkn2Gj1qqf02g1PUzDSDLNM9pffaLT5G4+vNtADdAA
1/9GuKy8CI0XQP1N9bRjdxsFnPq95Dt7IBANpIEIi3GhL7icRFvBagUqMnVN1jWT
+uUv2v526KWR0Q1tEZey03LF32fa9TgzV2aFre1HjGyiDxHDWea5LhLv3aM/Pyri
5YVb7ELdTXpc/Q/gxveVZtODxNXE076qt1Qp8Dk9chfbzn9zSRjXNrh7DyU1xPqk
9+S/cxg55CWYQBiC+wynbHOxoM9cuKJKNcWmrLVkaDV7vyqqmsommMC+cH58bBG6
/CubxN75locpSTW+PBWAy/bzWXkEHieAsZYrTIcX4vvU/CgXDLubp41MicjlX5tY
wUjU13P0idh62dmT3KxvHvIIFRGpUAPO9l2dee8v8gU=
`protect END_PROTECTED
