`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43uzEEHf10DfC76rBu9Bfv5SNrIqd0a72ehL3I4KZmuQ
KTDydJDjoGJYHeUum3JAx2zG2ohWlE64nM901SCtf0VYFsM56XzL5aNQ2J6GEhLp
rCga0AaSvJqhDG3TGp5tkaMxZWpEWLH2cxslJqizOtW7m3Hcnw/RU04Xpc3vCFTd
k169qYtvw2ab5PWnvffTxmLZ07vMm+Mc2V6Rvc3Z7hJLMgvVj6NFToVRjWQj6U0c
9c7p4gy9+h6d66Z5qpl1DzqYt2BMX/dShscDzrXgVOA=
`protect END_PROTECTED
