`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNyrhzdXd1niQz/CJaiqZpCmp+fyMqyEQvFmpn91w1Gb
a47+NEWTdXNDII3kHw/yGQFdyhR4zPt1K1ziAvEnjtA4vg2P/qj4SeNOAn95d1GQ
Xg20q7DAlShkSKbP4V700jI4OfLcsTXw3x/mHICXeD5RvKvCxudH2sClPtM0DEyA
7wU6BUGpd1690nXI0wjRmyCndpXf2tWIZsUJxMqqi/4TqifPSWCsBFBBq+6b5ru/
NMMOjwb0tGs0kJA5Xwrw6nisZpfwMw7mzu9Vh1waojuF7eQ2rfKcw/cvPemHNDLe
HS94kUyOtcQRdaqmGtSDBZq57NbFrGDg1fvi8Qi3zEqPMZA9ufkM8/viXyZRiIgW
O6OmFpn047vb8Du0DiWkrSlpowY49eQAr59trh2DrMsIx2yh9lwXDxKIX7JJwAqE
9Iy/IYCmDVKSuXt5X+Et6hsCP/gKpNLC8Ts7f2btkMBFKLlhZxKLYrptGaGf7LHe
Q7Rh30qS3/p6VJWhl83VbdVqq72BxxANjM93tOQoge7iBBCF114LmyQuhkfuSpIr
Eu2Ibf7i2A2Fw2gZKHnMEijGWMVvEiqDlsy/QAEtRmkYyebp6354vhYFGP8CoRXR
RUVQ8wwwxMlupX7Fy/MiUAmb3zO4RGCEHX206Z9Wm5wbJmPq4qu3Hy0ydXZLXuUK
TPpDVDtSww05S5sM4RXXT2O7Tvo18mzJt2KfW4Hxk4t1oitqGe521XtFTctG48fU
SBkHv7ruDy8O+qu3MnqtGAOuDM5Ka1wuYjbCUgUrf+vEm940By2e3QkfUsMQcndV
2PX2pTyGAon4dp99a1rDlRLAYC/IrmpbbCtNT7htWoc=
`protect END_PROTECTED
