`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL7Ib4MGmYpq1Dclw6rOwKCj3ekj1ehfampVfDfhA58Z
w5sbN+pH4FgPJl05NvsJOTEpJ+3OOEYg1AtNc83UKEi6vRRi6DAyun564moBMRmD
IbxaeXixgE+ZX0Um8EvMmG6FqkvxhNLd40nv9ULH66VlON0JhHSE9wjhFeLASc+v
231D+N+MzfyA/gjodM39UPieXxtpHd2DqxitPoeTxn3xew/TSfPrNYK0tR2kbn0C
XMGEPMZ0Ci6Ga5SPyEjG0svhCM2nhteZ0jinoc3+RSxXVbNURyMw02DlbLjKDbes
AL43KQ31T+8o04d8oH5nm+TZAgka9jkjH8nFpjBr+29mPUS8ALLs6DV3D3jO5r3H
`protect END_PROTECTED
