`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Vg7MbbcfROgalyduNEKoC0/Od3gUk3e4Ye50X63qNH17a8cPIYjAw02lc+H/gAoc
I+dXs3fKXx1tRn77mZFm6rWk3ndNc4kUtmxVNpjyKMFsOZkMJUMMvZQsuF8gYXnN
zMoMlTWn+5zA3R7QmTkyRD0JdkeRrI5xvCt/bDpJKynxbIRnzUq6/vjM++MHl4yG
YUmwrtzTHzuoi0ndSUlLUCGqcflRiyqoutJp7kB/CZ28n1RK670y7W83K3+XYLiI
ZIqA3YbxlIYsdFW2+DQOCP+p7HcaDlavLX5Glv0xItY=
`protect END_PROTECTED
