`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGYT0TvMXb1SNfBf+gYD17GUVVps2zFkcJ/5zCaPtMHL
l0xDP/eb664WUp1dhZWe26mPVCbiFhidIpzqfssXEa6z9k409unXllMI6DjZRMC1
2uKL+4A2pqojwy1Wbzfz9nA0sgF9MoENCTsjFZ6ypNm6ad3pr5Sa47gf0GvUI5Xv
NZ6OyjcSDtLrbL8U2jOXoNxCUMJ/c5cDCS8RT3eNTe7mAzo7hhrbBlyJFWSyW2c5
KcH0p14FBZLj7tjv+ccprNac5WAsEDpzlSjqlHRmBbvYIf6h++2EqhprIiFTSRPI
F8a153nqgSyR9OAcVkVkDlsHpmfRnz7uli6cKUie54zzsB/e/trjmrVALGlEZtf2
hVOwHzERSnCK2wjeu/uB+kBK3iCD8lVAAW5cqaz8EAF3gcZxxitXZfGHRhvQJZaF
Q7suYfcNfq38JT6JIBBDU5S9WqCdTHFM0tUAqmSR05QFvvRW4csN+iex4d0WWkyy
2QT0GltchRchSy/t8weXrBkeOZIbjcNqjKibGV0xwIj0aishY2JqUEbdNpEksodW
w+VcMJNvqy6SEh00pcNNM1y0Q/pAo9jq432ZpjdA6qE=
`protect END_PROTECTED
