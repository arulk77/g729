`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu477z3RxaXOjR7Pu8SuN5NuOyv8B/yfEp9F9b8yFYfwdW
INh77P1KqLsvqqMLrj7N+nKulZlW+r6ovKf8BR4lD8YlVG1VUomD/7sYD4p1t51s
MFjD7ORQ7dO/vHynkekZY/Fsw+4eicu0zssPhcIQIWXGMd4sJd6y7yA4j1xxOGYX
r1JiKmObQI+HgLfz9vGtALb8F/GoQOmPFT94oit40Rp20H6eoxlER+ix809s84i0
LeBeyXjZ/mnoNwTkmXP2F7kBwXKwuZXs5n/BD3jBon6SfK2dcUt0hy6UgLRJ3jCL
OS0mbRHWdV1hwDH0EWzkr4AF4a6FcC+cphwh7prqcy0WkZTIEptN0W/AZ4d7IYd5
33M7fK+B8GGdLuon1KLQi0BZXbFJTvJNtof5xNOBnXXKw9HnyyUKhTErlnBG9Ajq
0zo7i4LdIoy3V3qcBmiWFw==
`protect END_PROTECTED
