`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43tuSDK/p+uj/+cr+ygBTO+hsIZDTpYqzG70m5T8MTtf
2/oheVXnzjUgAorUqydKALcRxtDJ61m7TypOCqP/FslsccsZiTy2/OPoBYdvweaU
3H7o8MfCIpkd1vI9LbgI2QvAwVKiEg3vR39Zn4NxaAASmLkLkkQyfcvuAX/rWzre
meJDXfumplAJH/nTZQoK5QmCAEZneYYhPi8gR28izy6SSIX4weODLU3GjACkUt77
aF6AdaoDNR++Nv5sRQvkbnXT0h/o2hIlrDhyYDsaNCyoMxfv2nooC+Pny07Ai3rc
c7p+1M7IumeOuZeNZT7S7TqPwtR17MH5npXD7lfTvh9djh/anfHQTNHucyWz9IcF
McbU1JtDLJr6YDD9acgzvdlrPOX2NoiRX5WM7jdzZk70bnEv6Fq+ctRzL7llY+uv
oq9oc8NOEWX6WuOQC0SIH330s21/QNIzaghvlMSkMCUpglZOo1ak5HX8zvwpKTcG
`protect END_PROTECTED
