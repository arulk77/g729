`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu432Ix2cpGDAJK3FJkLM4sK0h3SaqbYKvgjy+Xr8xTmEI
suGEnqLwF6BmbnTwh3BdjGGHW4uAF1SIl+MS3QjqqpxEJBP7zYYJRN3AN4Bc2B2G
h2N6oAxSu91jWb/G+y4qdUFNzXzeOSw9PeKKtixzGi/RhL9FXUZN8jYP8idNZw2P
vjb9MoPBlbQ9u+rHSc/AQ23LI1rRAn7IpyG+ETwFlx1S2o74P7PriQA1KpTBawC2
jb6X8D91EZzBKBtLAWkjGOUNrVrCBCrSFNMszheV0yyCaf/MBYLUpRnAZ/A+88Md
xAygcTN122AKi1coL5N1EZ0neC7oXhQjg0xRb6bn2dL5CPrlSWqceDV8phARbaLd
4HyYrvW4vFzYjl2V+jnLJw==
`protect END_PROTECTED
