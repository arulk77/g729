`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDOBeSuef34tArGrK4IkhysZRqQHvFCtr00+FMI1t3hc
GP+PHuMberdEIw+szWzxMKWbxN+x29QdSF1wvcCE5XyFQpgIob9MCFCe4BgrX6R3
9ROo5nLwRVh7Gklopk3mXa+21SS7MMHadrhNrMFl4rkbxsM72xz9XeS51pPhEOdh
HEgzSluIC152z9eJvvX4ahmAxIbbQ6EZMGqquJ1NJc7UVocTuCw6TqVyn6FJas0l
SFJtYMYWBYZNQRNBMcMWL7MoszP6XJczXG7ypIAPS7oXoAxkI9vmagcxSzvbjGgF
HuJrO/iXTiQv/PpTq+dyMd8OQNKkxKkCuo8M1Dng6NaC0xW038epreXOsRZmivw6
`protect END_PROTECTED
