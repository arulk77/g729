`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNUPFrovvSYkBN8buaJ+UZGU7MrEjv0z0i+w/q5xWkEz
NcbtCZzXPHEx7zxzSvh5UMNixahWU93Ll/omMTHjv4wi/OxYfoQtEuIrl4HciFnz
EeaZvMpUuOaVHvLnVwSygMQFFMkXAm95VbUs8Z/bPr8CgTQlq/vwjyabPvNaxmcy
hdHmEdajDtN1IOl73yNcZZkqUlEEvQBBfaEP4SFlUjAbnpbvq7hpsVkXt0vWMHGK
`protect END_PROTECTED
