`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIAPa3ImYxFSz+V9sEIZQkczJiTpoxu7Wn3jzfmBGmdF
9iTeeFbkJjBdtjfT9Zr48+CejK7npfyEUrc11O9ACkoA5TF7s5xj9KatD5EORf4g
j0cIM7eofLuGLgQK/QO5hWIglngk+qNDdV+lxUVQvAd3tewvXNTy5JRE7sSvkrgf
xfLd+27MIQBBMNGHIFghuea/kuOvy8qOu3z+d9u6YUV4bGXuGMqFiprF0ORqSOeT
`protect END_PROTECTED
