`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aROGO1lTkB8qSCLuV8R93s3FWju3l5IOQ+HrQyrcI/kB
nwPohTrgVx8dJg1kSYg5vmI9NyQNCNeKS730N6XmbV7NYb9d7DQfOEfTF4xxdznC
vyk7D3B5XHlNE48oyGAjNqorJdTj22bbBdWouI/nHxfT41U8F4utZiR6k10+M2Yk
HFcTW61/8lGO9rr3TWPms8jNosBtvXusDer2L8xwBMxbiqshGf9vqQDg07HGftjS
hH1tJ+WkiztHDBD1FBLsPQS+dAEXJvbql01zrNdQF7Z1s+f96pqn8mJTRVlLUt9Z
iADwg/m37fTVx+wSM5bZRu8ObplaWE9IUpq8ts5AfFOua0Kczg1XrOqZnOyr9J1w
cuayQs5vMiTtq9EsAStszjiivoRnrjL3fHN8K+hQQwdwty9S+fKj5TO5gE4jh/Dk
W5iqheUpPsFtrR85HFjPP2OxF3fsxub5wZd/diHYpFTCeMJL0zREPq9ztYTYqBzB
f/+Q8tTCwSTppa45Z2MLzaGftni2BQkdBdvcWDHJyaAGU8UlSFTYnBWGHNYsqtFf
0UDJ+o+mH2Wc2PhZ1KEUGs59sm+WdKHTuFN1O2wKIu3lAswGoyeCzsb/lnjxUM3t
6dYdcu53xCqb1D2M1PTo8F4LGhoAf2BkJv0qQKZJzEkIyubIUPR4Q87ELQxGAxn/
9jkpSlI/bxQHbZUZDgCZgwCx6HE0loRXyK1l+Qxtz2cJfG2jjOf1CDVW6NiL507G
aPl3MhBZ22/EtAaSb4oo3+RtfPrjqyySinm8zMPFUakWy/n1r6c90pl1q61CzDds
8831p4/W1E9eEEZbJCEmAbUeXHqB5s+gdEaELrw2PTlEzrLTZROMUlB/tj/Ccb2A
VBlc2I0QewBXVWcoEHpZisAsoYBKI4BnsgUvQZ1xDouZAR6Kes0Uwt8UTGZu4Jaw
s9pMBaofXLK5YD24Jv5rkGpGx3thyTu7ve1GIbomNYHkg5hGDjAeUfs30e7pLaaK
Uxu4JbecIZuWJdDkKDkuNl9xPAjYe6Zi3KVbwrJPhBh1X51yu6d03sv3tYTQ6koB
qJyLanNAdhoUdpmH9Nk2l0NvoWImiq2I0uQAq6Pr0u33kUAZWkhQ+T6CJNlj8wVs
MQzkLQYbsoCybbkLe3MgAfVmflBXw/6eKYXTqrnMM+V5vpHo1wZxlxRNoK8XJoHu
i/gDkRZ2P3U2qGvl93RM4otrIw86rhVGxve3xTPKIQQf8ZD+cT/WgXx0sDartRXM
dtoCaEbpI+7hKQ9NGyjvhCqHhoNj+HQvnZFRhTtfDMKA6wlIxHo403OaQAqESpel
RSVidUXSV66AICBubl3LQj8yYD+YeQT2nm2PNQI+dpKVeO5/Ybdzp2JyV03o73LB
CRk037kHeYESNbZPCZXgz7P+FFFNnbWs1YU8CgqBMznAKw9c2QY+VFHA3+I76wZO
MU2U9y23JHR/gsgZxI1RxzShbrtgpkvyK0qjziRncmBkODLV7I4TcGWHZ9geQj6L
OI+31hxwB3hVFxkQmEmv1rdQBH4cqh1EFBif+ydAnFBJnHBOWvWViYdQXBwGsqN0
VpEO/hYII+AMIEbE9GDMBvlwWLrLrGAmb8Lmw76EawtlZHUrkAKd3hjBRm7WPUmt
yyIocMtKs/EQsjY6S1Nd+0RCHf4jdXVQdvp2avihDRVvhMaNABXUP8je9gMkZ6Y/
GgUrFBqRh2PAK7/0ZR2SPHyXKzu8hEqGICk/gDCbMYkih15+5a/3GsyUIEY8kyZS
25KNyFmGu38JHE6kSVQfL7woRyhfiWCTPIq6+VaWyrdyK+dlgfyJsbWE3FQuTnN/
+LcTWiaKJ1LaH1Hlzk9eReyr6rgOHDmMX/3ci87w9PTIM1jh6q5hzbVW9dv6aeH+
0Q67Nh7QV4EGe191GAzKJPr2xlLVtDTP+4SHrMm0ZxwZiSLy5W0t0H3g6xTaj9QR
TIy+Zly9ja/oflZBtr29C5lC5EoNryybFcmiUmKhAzYjdw6Ui0DGFIyn3WtAoaMU
alMg2iilgCRn6ovJJ9hUqEDp3r0JlR/+TaO186PKgaZ56CJw0RAVgJ7G0sMP8QoH
3YO06MlFdOF5Pa+we+YXFHXoTpAZ3tM5LuX1jJBEgx5ubA2it5t3Z/dfvZgM4iAt
vHv1siC8gWJicDnzHcv8C65C+pWAEOuafBoDTOvRkyCLd7Co858f7hMoiGouGORr
7vo3V3ZPjguXBjgM7KlYEPpp4l9BNWOCtW7nbrfilL5iBRKhuxftxp9IAbaTd8z5
QvFgk1S56rGJ4uJ5Rd2x4k72zOgsbDA8/5TSVApM7CArACPOQDJaaQjXuTUBoE61
o5jOSs4gE7RRjE7f/ibFpVzf7udgyd8IbmWDZYZTDWDRpaEJfxcKXqamhQ0T3PTV
zy1uLUkvo2JUsx3Ck2CMxhMWPCl4rgvuBFk7J96TDS9/ODPKm12WqUESCLEQwbX6
kB5MBBFSTFwda5hAWrkuZi4bwSnfyO+zx6u77zrEa4O1lEgqBfhqGyu4rIv1yWvJ
EbkPgwzmBg/0QWtzSv6+o4Eh7toYZ2aTcoI/CGg83HspPWBj8/uXFbNAoZDhIPgb
hkE4kDkFYQ4e4haxBcZFF11wLwpuPMh9S5VzyNiZ++f5Q3Aq1Cngj8UcYSWriwED
PchZyaXnjhiZFkj2ALFquDeO9uF5zsx4OYIcq14U7zgj4Sc34AQNQercgSSy0Rn7
+Rm2a+C0mzSSBKJnPyrCFQmTxw+dtMsYa7SYRYW4Jux1MVHqfygWsjwgEqjQp3iv
dL8EWIV3iqN6lQESoEprB9Ful2rCDPXlB8aTPmdVHQ3CilnDhV6tJnw/vqNukIQY
ffu4rZMPMqQz6ZZwATeashJHhzjRmLuqKt8qjDpx2mEEXs5AFn3b/eEtroSRzQ8R
6BXYJH9ah8k7F9+gxDauINoq4NcS5zCW/mV5FHigAMFl13oEggnW3z1HURsbAgXA
cDWfmQnpBzsepoOIStw1wku+OmQlmjtcgn85fUPuq0Qf1yMcM27dc4EFqdZEadTw
2lLdrFioVo4ZhjDb/vpOz4PIl/bA2gQ66xFCw5i1K9azxci8fjB7zzvYttrMeUtg
e7VColuq/1x8CLX2SGDpjALM7iSI/beqEg+0jqr9R2VGg6qMg10MfSp3IxS9s+BD
I/T5gIGewlzt1S7gJCkvNlCyhx0xcEIvr1hh9qDftItP8YCHuUICIquHUsDDAvLP
+8BSOapcfzRigW3EQQSAI72RQNN/4ofovf5HiGEMXv6dPUk0LQbsdPFHKHkeN+sz
zb44nyxEjBBvyvfSr/c8JaGpymBumUxTbgHRPQ4Zg1IJTY/A0LXKvxSFQwhWsejB
LyNjGpvBP7bEqFNBcmJQWKUOxSVjy0XuahVcNshwgkXmxuP5YhsRxZDdMIBwY074
gPW4bvStm7l6ZFVEagGr13czA0y32r4qAZJ7D6r52DxRE16IRMt4+AbTME3EnK2X
5xjnhMwvfhPcrX0qTIGeR8hHq52wz2Axb1ix9yFTstCe9J6PntNXCfzcD6vdIsrk
EV7WQAofgE3/SSssEVlDX9LmEpodheRhXzxUyZOZe7snWrf2WFx+raiR5oCm75w/
HT+N079uUQkgwq3m/SEp+0GwWWWTcM65VmbAeKX92LubGNzcVOZtoG6eeCGxKknx
VO1cY5Nmv/NyGoI6RCRPJ8ktcb1EluBb/U8XFbPto3cSJKZHL37XDmmtXRy2kzBh
Ozf45MoPJ02nmU9XQW2TFg9b/RmmDILucXbyamxCDuxgTkfOMT+PTi53UQxWGClm
OuXYc2oPRiqvIZcEc10U6C9ICC/JllTnhNfsv3pPkb8JbU6Q1+W7Hgx76IwgZGFS
GpeDzUrwf37RtE4rjRJLKUdSC9ELjYxEDkQFoR+ASCv3mJod34ubN8VSBe1BUQP8
sT7DKRTk4SfM6limsah18ZkezVIDhA1m5WBWrZBFdC/q1kMyjEkZ1jSSp3olEKxJ
FSc4DWV0i8LHNx2mb1LLMPubEl+HkokkZAGKHZE9sSpVT3sAAqHoshPGytPZlOpA
79kpQ+G1BKI4rIDE883B5r6KtHfz7E01HLiWi5dLXrc6FRTzehr1EykxeGnC8zhA
j4zr/Qls6o2nIjlwcZWOWrsovYS1XjOh+s7sK63+5tUzAGOha46gPdZCWWuRWOll
ydBvxYkvS9XdGAwj2/eZQbRxBRGnyJv0osk0W1srK4xOcS7Wd/qe6IORnqC9u7Qu
JNGdEX1IXD8d5QEqXU64E1VjNTOgA6g7H1i8SlRr1fGPOWb3oVdlaGE4bCE2Ahzw
YIfL5kloYwQmXjqBOnUGSGKOlpx3ZCAK6esAgAnvVnJwEVcqtuEp6CqE6kPDM1Qg
7mo3siYKj13Awp/b12/DtBZnEHkbcCURgroqSbMI9PBUhmlqMzw3pGbxuIcHiZSg
vFt7Gq3NpLeftIyZpzO2NpPh5fFWm3+60WnZu3xYo2gMTxhuYuujAT6k35yCCEOY
MtyE2peRrlzHeCaz9B6L6OscZkYYEQSxATUj+BmHz+db6cDC9zN8Zvnc4bi678PM
HfwBp+h8wEHOQcKwrb+Ezj7/yT1ugQdjoYHCqAHywSCIJRrFBuI0dyuA2hEoMF83
rbIYxIfFzG98Wzd6thStBk6mq07q6aDNP6VniQ8lV1HC7AoDEJK0fGQzPCzfBIcD
o0tAokU/qp6QLggych1CfiRGLB+UgnNCcVnprhWLkDfaITrfUXdjZYCqMA+M2Haz
soajwwA10FXI6XFjhG4O6YZgBQkVfDmEkuM8PwNwlmbrYvgZSHSz5L20Q88+Tb+H
zfnVHvGvr3SkC6GwTPHIRbA+oiXswkCZVAgbZ+zvARBme6IYcE1RRFd932MjjO9v
OBwNByOF37nR7jcFV+FRwl8DJUibFNjC/ZUn10p7XDaSVQTX0D2XHmN9YD1XBiFX
eUt7bGbxRu6Tgnzf7LcClaymkntfuCXeAJvUf7gndsybvBIT75ruSMzcZ2JDiYhT
A+wURdtJqfJPkGLJ1xE1eAEyWf23FIW5NawexXzN5dGLWJqP6jCDNiJboTUxLQGE
gjskhR71IqtQ3nfkgMsk2tdKcyeY4DuqrI/0kvdrXxwSLROk7+qYy8KYKrcTLlC0
MPCbCWa4OuzGTVlpxWUic8hzWo+q7vYRgecz0q9vEkHnRaxOelzGRQ6dKGNwUXdf
4lZFh0ib4TN1y1JUklv6hO6DGvmW9t9ygE9mwxWI8tLDY8MUxMiZ3ED2h4bg41qf
+AtrUpuYl4xU9A8nCbbiXQeuhUEXhExsllv4qavQMZqPAtwOmbw441/9/K0mCmwT
a+KeAmRzTYxmyxHxXlHw9Lr/SeKUUiWzqkbe9y1HYs3g6chaRMaXOTXPJbXFkorR
Nj8PX5h3b8EvTQT2Velgc3cS7XbUKxoWBCBm4YjzsPWV4rBzaRZSDzE0RuWn+zht
6n0MMfbyZguM0BY55DKD/nKczuZajqN72BlVmDct/SL1++NG875lxpIMBaJZpsS7
oaPW7G/Mnd+F/ZNa0oDiwRnaHBJtZ7z9cMzc1pzVmDMBEWCPOyU1knpGJxclyPqg
/Vqh8Yya6Ble38j51cBYcbXemY0aBh3TD306kNr+0thw2jXchZ39Ch/IJ3vNQdu4
NaQ7vfNS2GRtWPXNZCoEv3/fGk91j2xROFaLaxf7xGXCE3IC1gVT8QSUKdrQYhG1
ZbQ5Ts/YIzbLrbMh5qsSyaLcc6RlcK125xZLkBmU8ul76rMGhGZ2/Gwft7yCb63x
7WkFZtXJoEOPPHzIQ3CWWR0n/CKAZX0Zhd7qzJ4/hmnOFcE0cyjs+TmcOlIiXGrs
j8xk3/V9gG6ZYrngHdVesfF5349cpsmDRHitvUUaXQVcyfa/CdGCXpHBf32OPtbR
YRBamChEt4YQCOFRosCUAuriEM6jYDZNcCAxjFQKzi0lEwvM0oJNHTuuLOhMXUWl
QuNG66KvI/CaQMZIysmVoUeDhnPd0UfXNN3GS5JxVD4ZH6umDFbVrgPLNce/gkcW
MUJ47722TZrI6FnoXgWg558DI9CuLS019USwTCcspcbOLsjmSMJB573gMVsNGF2O
knCm5OatH7RbU9vP5R5hggWJpX+DA9U/4ZguMvtSug5eKuENKxNzGS/gc/NG+cM1
kf5IfXG2xfiZ+31alx73qpzy1OtlQNGQkTc+2NOaGB04hDbTSOcL0npK7Yo0dTJZ
7eUF84mBbSftXmxy94PHmNjsrNmm1hlANSbHvqUwwAhEfcpZR/wgHNeCXkClzyTO
VKHopvh0ReHTsASt9IiCx4P3KR3oAy+Om9XY+SJS9TFcPZ6hbFzKlAee6FOot7oG
WHnCq68vVow5Qddp/tJMpjFdHOSLGjRdAGecl2QNRH5KYsMsdjijxIAtK04YSo6n
wd42lQD+MwFOsoKFnRwUu3TVREsBQ5wJM+XgsuA9IX10htGSWqKf9cii6i7HYSSl
sUM1LNRW+cvzPpcxsAHIJE8cXRdj0sc/54zXgv6subI9EFQczswvChSmq2UxwV7l
rUjjA2MKgq1Yjt9atv6IyI2TknL4+oa7wxm0R5biCeGGSXlE9hBT79IQl/JP0osl
ska1Og/0Cz/ApPdkiGKn2nwd0b0WxOl3jCPZ0M1kjr2OyD3rQDpmIc/5MM4i81s/
CBj/eKe6aruLfsFMviGQPGePJDhpcVyy7t8g4tbWPLQDoiNXH66nAVYmlYyPQE59
BFYa97q/fpHaVLGH4Iyv8mOYSKjPEd6q89CV1qEu2KjEuR1fTtlzA1JaXzwCKxPP
txBTCZSGBx4qEXLsRYomFpJmbIH4WewnTvMMjciP6EBwVzNwLXmKwM+aQl0PnGla
zF06BD3k3/yIVVHyUm64rCWnV30EGJM9Cn0QgeHp1MrxkUId957b8QqvnW1cjc6S
dB6GIsza6X4urwdQOnNdfXziXSzGk6qjS3rkDLKQUkv+8VNbm5730IKUODSA9GJ4
P/fHPV1jaPmsErw7I0MQnLmkDPeR72ogPTmLIcp7n0lUOJWPJzQ7ziVyIpa5U+ah
VlVWKw1VMwKwvjs+w/7DS22nhiyRtoCwPTpEvlp6vv6ZoaZTBPk5Jdj8O+MhEVop
GyklPuXcSDZp6Xcr/3Ackr0qgN9ADZ+PFFCQ+EWFkbhBmiYZ/jDUiH+xZL528kRo
7kqEaFQW0X3JKFYSKmShnvV5t3c19dwXTmjZK0oiucyg++tDEIGo96fi+7yo4sgn
bxfC+Eajn4O9uFwb75hJzJKLnbGFEZ1x6CnPMimXepduN+xt+CWrMFB52/4I3Now
ZTrf8ODgDIQzBLEE6PlxbPxqGQee30k+WIJgXZnNCSnxxrkK2xhiOPuI0HtMFgFG
yqvyct7Qx4dSKD+m61uTOgIy2Mzl+tg1YqP3/CEaz+9Q0aDgIwp+wp13O5w+/lPF
7b+mMzY/rnP2W43WRgtP2vivD7GlbKHMtKF5WHd7Sp370h2rG3XnP29r9OsCbmnc
I7Rsom8fnSV5wgX64F8QhWe8c/v6pOZaTpi315CxjfhXPF70o0klz8gVmYtRi9Ej
xcQ0svJjKLUmVo27oCZvHZJNCJNpyfwxaYNC6JHSiHCBblwk+37CENNSbTzzimW3
XmXNG/7ANIWwWYeIQuNj6tUkFLU2mts7sm1m9+Yrb+3sY4aORk3MSWL5BornZydb
Pu8wSUxfUaXvE31jUAf66xVk++BesL6+5DZrO5W+LUOCXhfwZAgtxFxMT0AEaZrS
IrnvqDWw3zpnIW+ejiWvwjQMtgf4k60grLiByPF8hKjUTXeuT1vM723+mDXsF2Dv
i7LaEYUDcsuHtLdoKf/vxbqN5jMZU9rVh1j8OzK+5cDP0emOgDnb5qcx9flvLD5l
0VfcyapNO/SbHIZxkPP2BvM/R2BbLJjnw4lIjiwo/SIcT8/Hn7H6Go6dU35W/FCD
Efztu8kXnD48hu3L0OOKJ7ie+k2+CvfnVwlBY/B5+Qgt97syWUCyLWiawxBFRlXi
lqUIy1FQBLPiDU2NTZTpcZ5guZMPQY8qoPRFE1Az7yOn1aih+aa7VOPkSrlEma5N
4cp0hQ+1yr7oztiFub8uRcYPxOSJ7mFYfOHGguzODwysiaZ1RI1myo6kFXG+IdCV
m/pqHrxOeegwJtzbBXvg/sjgIvfUcLKXw7/OQvvxGhJtMtojq1cCxKzsB+0kC4c1
qZgl4u4vLdTB4MSArl1AGwVFQjrcemtgJUq6YWhUOiXa3wt8sDRV4Mv4TfMHFPHu
Sgx8ehyWl2d4wVzkou4U5AL9267o0SsXMo1smFyEHeXVtfXMHfvCA0E2D6yYiwO6
srwo78amrbz5tRJYb5N8DSX1U+40RTMRXqzLZhxT2PCFy2GQPVg421gbUQb14xUN
KODsz9mcNdbskUpzmNnaZ8BZfHbbPjbIVPDjxKJ+CTh01o98nlWXYzjXSJAJMrLN
nfiEauBVpxaUmK0Tlx5O8ZIhgNZ8Tb0LhABuTttLOQGI3i1wzp9aHF3KPcuvpwGm
yZPOR1DIcgYLyCSXi59TiK5LBGnct4NpLtrlGH4qqEBZ3BDLMrZuFuaIuBox1Gdf
ayh8ak1rNS8yTidQIAyPv6D9vtluqMaGW1XNTJIO1yNzB/nO4Z+6HtWFPdTJCO8D
2R4pPAj5WP+yIqEEZnlpph/CCKFsML1V9+xNYL/viCPJJ4OGbSWzmRH42CTs/Cgf
SHG7JDTAVwKTJ+qGRNpXoK+wllsAN69QtZ3KImO4dMyfnXjsegaw98CKFVN2QFcT
49SVa2TENNioaLXFGRI2JPeUhUMYc1iwhYG6KsK3q+XIg4JGYHc1GI4f9pVXxseV
v2Ya1KWF1eI6zkKjnJ267oKJtfaHft1HxD8YddE/dTOmrKRvrzQwUj1nF1CZmwbk
zm/YNZ8tciu8IidAlVuGPlsw/meBkjvwUii9stOC/12blTBytQNZu8J+3Q7TFqWq
2UtvPQi21OJbG7E2YNn6dJcAR1H59PxJlvI1u+IuYWGQZsl3gPbE3NmGP9YV5Oe2
ksNATtt3qGAHWZyq0K/WNtiXB/xMWb0PUR+wePbv/F+zNw1sXWn7ZNy/2EwE4jxg
mtAJmwzguefM4mU4afNd6QXbMfiAGH2srOvtSzME9P37Wzupp1Tel/Od2eXGMVX5
nnwkHhuehdQHL916eP77SgJ5HMe4NmpNMR+FKXUg2J31u2giQkaoRvA4XAmRW5Ak
5tUPtfTUyTXMCJVJWhJnYwKVjlZGApeLlFSQJrQNgykb3mKDb0vi0SqwzqlwEPpb
xoUDeeHPyu0E58yym0w9i8+aqhzX6/U+I0+wNhexngQgWsr0qPAK4oKm8pOq93tN
7DbUv651DrW3PX+2NzUI4L3i0OOcZ4l9toNGf4Yfuua5eMZpjU6NGYo/0JQbDZUj
iUc2viuYO8iR3fHNRIoD+EXb9eoaP+0+2pVGmh/8nAJorVbh3oPkiUpVrHqvHRBX
vEzBoA8WpX46tjcWLPMJdhv0uvH5kG3sK6k7onTJNuzTYnzJLU7PvLDRS2VEp1A+
465iibUOtgcAymfzD4czh5kJI7oJyplAtvwRGyH7sYwya6a1jtVhkSlQlPqJgkTy
0KJS+ZaLCW+BX125OsIy3wHwRXIw78qgwBiqIQXXx/XRti5o5DS7vKi3xgXQQPJA
Tp1vmK7Dul6lIp2nA3Rs+5w94FQINM6X4D5aImsbg851MTdtikQ/Js5mYAmqe+qV
CxfthMC72doF7LZEnYoUMwKCrtXL7dbzbmILDWtBKovjgfFE+PsvPZk1+KRvmZ/P
M9wx083TGvUQOZwAEJYFysAtpXNj3CxZqhL7w1zUl6QdyY2iaNr+8AJAc7Op43sm
4HwseJfJIUbF3tcj2oMjy0wCvNnVTPuxuJ4QwqLYRvyOg9ugcyvvgypk+XAtGLWY
EqkvHpfqrJSCMQsCGUK0nhFIl4nooTeYGNm+zU7/NRDAInVb99UdShlJDcKysA1y
qqj/n8qWh+diiEXPSD6+qX2tOUJ9o04ZXwB0GH6T/rDBLcTuTLc0EzLcT4kLtCWB
72naLjva4ZpcZVvSXG7nTK9EpOFrzJQD8oXnfkE9mBF+TmbWdaHSSiRaaX4amaZF
QAAEuoPDq91V99VQzvlJeLx/DkLcKgSDRd6ICBHeNBqruM26wYqgnLlDQiXYkRL6
kohuwjSCY+jISxVK+xlFpu2TFFFO4CxXqGC40scDUAwOa8eTYfYjjv6S+k/p1BAT
gE1UBRJnGSHnd/NY3d04Y3xWDYLgjQAQcSjCEeqppvqXjdl4/1SQrdfjh6Hl7qRK
Pm4c3byTXWaJE3yqmaZVfOi1x7KZAGDBbK2v/BwglYsqI/lqoUw59tSjHU3LKrJk
8l1LjmJvLn/XHDj8m+MSM+o7Pi/SFU1+7AEkQwecCB2uUfJ8seNzb/2NWB6PixZy
zKCi9CN1wAlAYYx9RVJIDXkG1UbuMlYU+rr8MXwBiTO31VdjQbhDozGwdiSg48Jb
R95GY6Q8xEVsrF7vthJcGNjQKX8YuJ+cJvDYajvH/vIQ1R+ovu470SmmjX8KytZa
Gbl4JdLHvxi+spr0/pu9kDHodrkDSYIAaRWVzLvswzJc7Q17GVCHJ2joAm+SEGC9
7VG/FyZwwernCpRZsJbvAJTo6qlxf62JwwL2AxN2Y7Vxc1uTB1VqSrpSoKvPuNmD
/LzD/w83WawHjdVcOrMDPxICUdUtXGk3LJyzEqLuOzCCpeZOS5Q/uj6yZlAZ23lZ
eTn/o/AlwHdHm04u2PzQJxZ1UtY0lZn7dAKR0Xjlk1XwT1CgOEDXCff3+/X14t9y
IoxoOrFoX2yD4H1iSJqCv1tOWMP2swoJkAzriqbGHLmQzlMrCTCjaN9cVh9DiK7P
mkA/LSW90GVXbJI8gyey4gxpEX6Mrq5ADsoTPq8RNnDPfHDCb1XJsown2x1qwDkx
quHAsKqxBU5gC5qVPC78FF37o7U68xle8qcAliWcXRyE6xtha7eFSNwv5utmhjVF
8MroIoJ05u2hyPPeFkZvfEf6l1bcojkmfit34QPkzYTSJdK61xpNNCzI59P1plio
Y8e4QTYcl7kmdlF4WA4OcyGnHnLROUYv2pDzJDVe4gw9kXzkk0jfEALDPBiSESXK
QsO+3Nznqy3cjzzmN0jtQqN/1iBfToANjpsrCUu/I7wH0bxNLymahCHrjnHB2sct
GVSBGQ3xRfhZdFMjynvBPSBQQ9HHx7lodD0xhuWAJr/t8Eu1pn9mh1yBuo0Dn1E4
KXETo+DTkflN3HUDQtDhLl0ka/0cWDuWEKicTK5LrFjspvMwqIz9lgFxpMCxtfgO
D1DG9m1pcqqlrcm1t4OnzJ+EkLwp2j7pdPyGwp2feDigPqNyMOcvGnoiVtQDHt4P
SA0PrrDyoibqULUBsXIxkxxvHv6gJrBGD7o03o6BPwrqCrwqWbQNmmluAJpzO6UQ
sTEuTBqxktT1T0CpnTMj/4CTiB4zU5pYg5d9XsGQP0/f4BYykdyWlbpP4Jo9dh/O
iu96omgKgHH7iCvpqwJ8At1HHp4ypjRIkmy7wUuksY5JbODwF5b6JQTqdIA0DbFg
RjgKLoWBnviH3zYA+S1KdEkZg9JAlszD2th7s4Nv3wspzsMr7CDdl3MxseY1U0lK
jjvzXp+vDIzCmluxDh58mCkp39+HtDJIobObBGKtn3aLdWBUogCi05m+2gFpq1fu
zB/pdjBENoy1anGeEB8nmpgZWA2HF4EBrSaS4R9e1YPo9BwQXNj6gGkalxZqb5A3
Yi77DWmCAdA3jI3y6Ps9K82b7WJzYN5IUnl0YiOI+T5oKXDSEhAZfdfsIy1ujAXY
yotfesGLkbpOzL8CjJUqZqLiQBxOXLOKzfy4ILhEwXWU7xMFZDLrLR4+jy/Uex2Z
WUXQ/AOIHOfuj9KyNgh2ckomc81RVQXOK8JBNAcrNxMI1wbGR4WAmyHW2/R8Ozai
lIO/eykzDO8JXBg6yp/3HZ8NgAdHAEtnMXwHUjqAhtNFwjwPPzkkCaTIywRdDr/3
6p89MzLDGzN9i1rSaXN/ScZCus5HMQsaxMxTrFCWC+fHFN3E15PqS+bYinVpcypu
Ohd3JYQxDyk28/F0blHeLlfjvkXTtoJvNE2IOEL3/FFq8EM+NmJ8ScT0k9sBeNRq
g26JUgWQ5fbPJ3h0CsDG0mAx+/4AunEt3tl8dpMKIxFtSjHpBLNKSwwirCitwDAE
Z7Nkp+kkH6GfEzVwBL4+7fJCgBo9yS0JttV27TKsKYHiCSedpo3wtzrVq2bjHWkN
t9mF+SzqVZVjwKkDv7wVp0D+8RgE7kq4/sK9on0vfxeBtgnONJHxPcANwcqx4mxy
3Y1gTGYaUKNcYsvmzUSVZ58MbgAJDhZtMYEPA+tk09RPIpbR/kOQ51tKOUJTcezy
j6SFm2EJswnHoUbN2WlVfwMgR82/bsy2BiFGcYpV9dkOyQlPyj92dzEH2ke+2O9e
Ys1iWtC2qie8ec0t9LdeNyq2UjfWraaJ3mCEDd8wo/JT++/x8hi5Ihr8JDEn47Oh
H6es3MX4qq3ddu2gNOdJ3hDOt+fAErqcTxoSDyailo9A+IxcikUS7QJkI8FEIjXk
9OrJAAAA2mcoUGv2XBwRce5adu469IrVecksPAo6VvwzwiENZR0+ffGaJUNr4j1y
2bP9Ks/QMqcbfnlJjpN9X+OVmeDpiXZHBw2XuivH+cdJdoSW5O0Rc/YFkoBHTmql
JI0sta7XF7hZEyxYf2AaMue+2R/5I7baI+nJ0QbbyI7rlwI2bSc6+UngvSRUEmVc
oQN0IH9oGM+s8wp97fbT45gS38WD2FYCbljnwLmTN98UTkasFs3knwnAojmJoxF1
uOCwrVQduIplcsNBBNVdvwInA1n+xrxM6Bvj3QIWlEUTU8LeRKOlXZ4sgCQ+bEUJ
RmeBJwKg+WwJGNrxAW/PogaqBRsFfwx+FZzvnF1BoEl+TtqB/+5ORDqyzP4AVLhA
1/0GyyxZXZTq4JEt3M3KC2XDu9iOz6oMs3Aokc+olPZGl1+dwTS8lXbfhPp0TBxQ
cgSW/vrucgZ1DmP3f7x1lowH46EllPcfdgpdwPjXrM66oGKXvANTHbh0jfiI5ttE
zT+XhuH7ozWUykzStpDpk3MH+MmMSoR6GWXgMTkVV/p5r6M4eHOBC46f+kzws1e9
RittaLdPCa1VaN2fnh8ArNXsom9GSjkM70xJ5crcRvEyrf0a78uILjv4s0yDWfEU
FBM280TpCAvDR+dAgIoZoqOnN9M134srX6yy0Bd/+w6hJskXZ59dHeEdYQ/OrseD
IzoojRmOI22mlqIaze4QGeq++9fpDH+QfdbGl09FvMC4yqcnFDXDTiY+j49p12aU
QXx1c4YGmh3l7eLQDCUGIfSwjXJEl9Owv6mNMYVPxYPV3FuZoG7/QscuVs7j6NUH
ZXAI2SAVzXF3subk2bdGnfq9KlfLzAHxhaolDTFClfNBvwEpBKCI/IbWwYpAeoTP
Ks3A2+S7fv/JUm+LK17iNEN0l1NtujzqG/9K1MgNUZUMo31P+ffTA+TjwayfnVFP
9cVBXaWXLQiQbdS/JqD7t8vapaEdJ6C1Z2hZXZwG/d1vTtg3mNx4Try78cghf1G7
vMTPEiZS9n3zbLeUo+TVxhnp8UWY8m8cnwTTWuWVy1tSGiEVIblIAQexeCdj0uwR
G8ws85k1q6yCh9w0DxtqAGIbk2DA4MMumR8+bI2WuXx5OWroKoQolYHNPucRIViu
hTBTIpRUSW41jatpa7LfZUmjj4tDllL+PZTCuqy4if4K79x8jD9X4KPWrk5rs6Q0
txq2vZ7u3YOFIM9+Q1wwJrppMISZcrWxK0PlYR/BMdSb5WjD4JRhw6ArTisNFJxx
s0CdowYqx3pT8ocs6FjyKLiR2PZQivJepWEaQNq44SSMU+u2cnJDWLnbJAxL5gKU
Ll5Z/iHbb7NfzmEPjUh3R4mwNES4q2jzbKo6km85kLRCgi4W65qNzvqOqz0gBsq9
RRBHNRx2A76wNdWc7W/Id6LeqODJzhfTzpWCcax78/egbpbVQUH8PEqw13qLSbNu
uYOQRBjwUY/CClThS9OMC1AiCRfIclrhF+LddlcfX8R0dRoc6DM196mkboTfEnGT
isOkbsnPMi3PR4WFTkCHpDelWbzDpAh0X6Q77D8U5D1hTPIjArUVMXnZ6lm3WzeB
mob88NSn4fdJ2oMY7BQepPLF/fiwualrrOIVKJteJc97JpkQiqvKaT7lEbqABc9Y
qA+Pjl/TI0W+ih4GGvQ/74whzCFls9E8sOzg1E2e6DzpjYebk3U5uNL3ttVucw3D
ilaCSRHgDIzdA9LlnOBpf6BOIS6zATf7YbiS7GWXqnc3We9eDFndbTSF9BlLUf3X
LKQ2yV3aOx+Niy1v158wRjN0wDxgMKQlK0LJiTpRn9wqhC1y9Ts+nu1yIi6GveBo
Cw2JeMMaD4RVlEZz69e7dflCcXDdfgpGpPmju5yoNKsU/3slu9G0HJ6bSeFZkz5q
Lb7JMeP99MB19AUXRxQVAOusgUOUOZhyxUDjvR6+dzEY+Ydbc2jdlNcrVTNCRP7n
xY8A/9CFUtsoMvXAvdpLsdVc5r5maVb9AefuHqd1F32vOt3iMc+sHm2msgzekymm
PNgWzMVSdqx3HuLuZkYo1Zh0KmswvmnDVT5zzJHXLPDZZZluqZaYg5MCEFj6tMnU
LmTo4VhB6JnSuEjKD30VaiehKTvIoFIjuWcYQFXPH3Zmd9HMJnnxKfOpoB+jXjUg
t4Uojt2xCI/QGjK1IT58XPXzgNWfg5SzKjKBabbyl51nAsEydeoXR0zgNOysqTm1
rrO9RnLfqZZttnkpE1chPnVau0fsItXMTy77Am+8022TvpUqMRfCzpvfrFz1biWZ
Us8ZCtii8Ku2zTGqSs8y6yC0l0QORrMPoYC8zoiM2clAqxzziUXp5ZvCV2hWtyAm
/hD+jOd/PvAF3fyK/Nt+tE5WYSQucwwiouyVjcruqqOyZgRkEFBedqARs2J3DUqW
wqoqSXufmuSXbPURMAdmKPoOduiEE4/BRg0cDJpzgXiMTrSDS/5hAcuYjAb9G5Nr
w/G9fCZKriUR8Oaauw+Lmnkjxm84gVRFoCf3vh1qJTGspdWi29+Qq0s1+Zpcux0P
2+VR249o6a5aZIYTI5D4iuaCzjJ/GDbMlotkZ1fuHNGJ0qvk6hsRU1/Tu8v3HV/t
AlZwmXStjgg6X+HrG9fQJi7m6c1SAKtIKrKwNfdzg2+rBsr6O7ZxqCWgmeW1LgmQ
B77uibhdWgVtt6Xj/VHRiUtEvwkK4+H/kmM9TzADuTZBHVtcjQIyBzSrcQE4ru/6
uxGVcvNZU/h8XBeVnb1l9/jv4v0BUzx+iZURO7P4+g9Poj8UZpAzfBVTyksk2kLa
s+h0I3G5WJI0PabkhnllvYn3ldNpdtOOQEJsMSvj+F67St4RO19IGlFWR1Kl5rZk
LpS24Y0ocG1hqD5bLn5pyxkXKE09F4fCALIU4OHnmGidh4YgwAfFMpUVqII8PGjW
Ee0DpC5jqx/Y0YFfRBev8V/VNN3lOQt6qxtyaPabUbs+YTLKdh97YlghPp09R1dP
qt4xCfYCeF7F+0k9u0zvDEg12oGfduS4rk1OGCDho1HUhc2fENG6HDCkcpgIFhgQ
G2NjDfv4tzHdgARXPOoSlJDZlw4ehwUgCrkQxqHkTy69rtOKMo417KlWE7z7rROy
Yc2ElpeVy6lTHLZUz5lD6iMHi8zl1pF6LTmlmYxgM/jtTJ2Pc2i8Ue6Q9fpJ7m+Z
u2KOgOGhrK/VRaGnzIZ/NNtV97FRZ+/98EBKMQfUAQIZONpxR8bYfq0MmfWrU66X
2RzCf6LkKzgt9KmYINl2vljOSGL9txo7J7W3mdqa2/trEbmeMh2zBRpsiF6X7atb
G+x/IxD/RlsxfLdWLa7IPWYIGaIhTvYg6t0S6rwfraGTrkVOvmLOxc+S6dHmSJ4Q
abInbq3CLwG6B2FQIjRt91WaxrsCJ8BAz7jGsoayUwN83lkgFmctqltRDXO2CIoq
mRy/EJmUw8dDFv76bLBwGqR9csDYhtJhnEZKUwbNxHRQ6aFBJ7g5rx+4syQCtAf/
YtQnKwHWICmq+M94fPtS/x6fR702mJaBbXUtgk2gmqM74mXxRXoJQR1iqSemkk8W
ydIm1bSccae9S+Xwoj+INswaSGmZ3QQgkSGMMSDDcaiJMfp9IINa1NdTI7D9YZwH
xCrlDtiVCFZ3kru7im69FY00+muWwDbwcHDR+zcs8HbjGjLUbFexjKSUcRZO5i0F
Rk7OOO/Dx1uWfVTPUUKfYb+ijA9xH+B8Jrrc2H77zvLnhSuhK6W1wI+bBvlWnG/D
+mMtltzMkx9LjOBcTfCAwT0CgFb7LYm3rCiCXZD5nqAiSut5XWe50+Z16rFHj1wd
t4IM6TSeNOHTztxD3ixSbkNU0QFfNER93sZCRW8nRy7h+oZh4NBXoajefOtKZbwE
6eFnVIcqs6hjUXwQ2nzfn1ajlaVU8grJYLGJskvjQorIPRovdPcacC7thb7aCONv
xs2lj1z5DdSG2z4AGBeOq2dW9SEaoIiA2woIBTSYX9H2auZDQSoZMWs674KlSSbe
sAAF78ho0RnZs9FMlvAzuVmMOr+SeX+BJh3G2dMwn1S/o8pyXPQynPZVyy0cLSNC
7ZsqYRDxWun5wH1ZtUkiZzE/xB65JUGLeOYGihzsXQZzkZ0Z1NT0Wh21lOyTUOVZ
T449sGWbptqLruyZ/9tFOHMWvyZBcKej5oWOYtoPTBp7gNBV9TpMd9T/7nSLL2q1
rYYFocJunC9LzCCDRwgskjNxUwfTO+7GkOAmhOxwHyI20LXMG+ZZcgZscGme4cRj
xUUdqhPL0IBBgGEEYa+1rHeCLgpDawi632BjbzQDNKyDz/med2+VYXTks8M3DJ1a
22Vdd2+XcTPk/chuMkkS82R42bZx3PO8cUUTCbI8WsfePOPb2OcoQE40JDX5Vvoe
FMdaDkeUW25Uh7TyyJ3e1S3vlaEAC4nBirLJ08dBQ+rn8frncVxvyEzuoebiDtTD
xGF+TF2GIwP+HdvdDI7S5F8M5CnMmPDp3NZSGErQr+0p2HX0ctdqV4/qQExeK11Z
fHRc4QdGCoAAaPQn467rksj9DmZtQvzYdsYISLRXpHvQvwLX3426uxzG/6kUsqKA
KGeZZKaNNs72iPiNXkO2jUJjTxCJG4q6KLprwOPIA6C/jau2q6FhoGb3V/eVuEF0
QCBaKwwQp/kSx3saXQPs6lc7jLhE6xzgXqeOSawWUwIjYzo0cZRtK0p9wUrbWQD6
e8O/NsHXdaqBElYmYNaRTV/+Bg+hOSxNOfYk7CqQgjuAGeOqJ5NbIFRzyEg18pQV
0HiYleqSrAIL7/JNDMsGpzN0aDMgnmorwgbi0eLYzQARPlOrREKBqtBRbR/EjS6p
jbracVIgPtY27M9DtyS1s9sbWOrR86QEcwzc9OxKcPiI5hySmKLw8FxQFTkUxJwv
lcWiAs83AJjwfiMcaoWTewgNCyE89DnvmHhK3IDMuq1SjJ7pWi9WBSNIsYfrIYkS
zQ00zGhf2K0YI/YJcpgeTUswN0al6NkzdfB+GbcpiFpdKd5TPGWpgdEOYRYcMRut
BHoJYF4/GiegYfTlMNqtcv0RrmbutDelLi4xw+9CJaA6QO+LZHk/nzDLKeKsyA0D
TyGYJn6QRuya6O8io20yn1UHZ67lRbPNcfWhhPzF/RA/yJE/k/zNh+aoRdjyizCP
jbaCG/zkbmPBzUSmUo22VyvIg7XULLTGjRn0/6d4V2vsgrYbha0nZZ4rnKFKoI3j
x9ppRmnqpjRnMDhZHLJvOCL55nu2QQ84Iaet6uYVO8EgtleZWuZngrwtGYHpSA0d
EwTAu9kjuhfDSTEyIpM2s2Kgc1Hzm8Bz2euujI6gXg2qUz39rvttC2pxkcNFRgON
uBTdbpsblaB+lkT3mrbQtAPKLupsvMiOAw3/Ya98bGVJGfKjeRY7ruXPOYd5TfpM
+vezwdIr91eZn2XdRiyWp/jgM6+YX75+++Uks7um/TxlvsCujjjMxiXe2HSAk97/
R7ZUe4/ufklCfR40INcAb3zPYL+BOeuFgcYSuDdcM0XwRL8NaoypeRf/gMPd7ILb
WRtqE2dj9cCGicnXHg059fGpuAJ3rkhwqZrzlw3cishajZmUFSl2PZj0n77/1F+U
z1T+lGhOIWF/OaE7WTrxxTmfRrZV9p0q7+/vs39CqD46Std9z9fphqLjneZxGvYp
SxVmSiA8XNPf/jfPkxox731Y+PCEci9PLTrDkuS98898Udfx8zuwsd0w1KhQlYkR
hss1zh+D1geDJOLw6r1F3tvfT3M1W+O9wxrnEAK6iBEJZdUOZ75LEsKm3VN5djNw
CX1GKn5T0+PU4P7p1nUP66fNrPRykMbWeVplD0+6DGqNu2YpTRDThOkZKcea5deH
2HeZvUzHsLJn2jSgNCFjzpDGCPgbDIgmdYIWiz8QUAZl26c8JvMGv5IE+7kNdHl+
AYJDlZSOMyYB/hvILnD0mNLeEf3Jknjy+Gj5MvpzU/bO2AWVBpB1qItONw7mF2J9
itAi9KwKQiLVfvkJBJVQfZIEWfTL9hGz2sBRHcaFYNymj7RrDCpjmb73qvjMmKpN
MK866Rayd+XtiRWuj+ngUIAJviaPyN1tIFMTH6ImLPYC2wD0sq9bs3pjmQd9tdua
jpBRIZSoI4kznLg4gRCgyymU+Uhi25N5FedrDHzixFmplKTDSPqds00j6VwvxxA0
XjxhWvBfYpF4bF52Zei7Cxhtt6Q+R8zDn2v+qFilQ8Mf/2HM8g2FsuzCCpDmlgrV
fjp+MmZKMiLYHyFCgQ7vPoq+QUsCwe55H9cl3u99pLq5G/aTm4y8ZVsplb6lXYqk
ZyDYvoaMf7Kvo93up0zeEwoCQ33RP7WY25I/QDLD16UvcJo33ST84aHz+ukbp2tH
GDDd4CJcCgmRZoWyI1cSxIKcdStzFYuyPbDIchrk4YB0IdYwrJxsaOyXJB1TCsjT
7zmeiTr/XvrZPT/1V08Yqn6dMEJULclH0OR3WGX63tW9UNULXhtN8hqsZVZ2KImy
cqks/5HXmq+vAw9+q+uJrUcOKvHaO5iwXP2Hc9rajXsoUVMo/fRwbj3m80mtsySq
mkaPbd+Z844iQKj+V0CEqJVPi/0B1ntZ5sSAyylHGa/ukMCgkLRN9ylGBQRUSX2b
JqMQKryJVna2Dl6an6DvKmymRGOvjn1J+qBmQ3CX2YzO7ixDnnwKhgPbMdCuVENc
yL2wGkxgzTllEMZ/ArZBQYpST+pzEpGVxojD9pkiQMGG2wavt9SN7twXNwFWvUX8
bF5fkNxtXKxp5yRNBlFjIniTtp/a6WZWdJ8DbStQq3rCGiMeXzSEH/zFNZLkrvtf
GAck5mjNKzKGgi2L6aSSwlc9TyXK6F/EsdY5o86ND8NNT7B7NIOHkOArCXi8wbjg
zGXZsb5qeu/YLoKAyZ4jyIdKbGeH+8nzzaTS26ql1ukYlOaBK08ZhdCsaNvkGObS
cK2QOLAcopC8i1hh+Nf6Ro6CYn65WXwtH83SI/yDjGMcmnzUUCjJ2RlgUQfaamuy
lyKWbgzT6kBbK/tHW2T8WuEUxwqWsziu4y7zSJeocDIEZvjjUtz40Na26EWk0Q1w
9Gfmm7vc3PQ6dynCHymXpsHOTZbrvf6AsESexsoIQwWHj0Xqsin7sfPTsZOy0N2w
88fvirzWwkvmmaGWV8gOTvsVF9/9AwQzHLuO4PiMt/U1IhWhtJZ8VItphFL99YWx
hp2idnQXkzOUX3CQ982focrt/g694ggPkkysktiiiyK/N4QEakqISzqp+sFUUVUT
hP5XRSUIhq8hqYBdb9/H5lcbbGgQTDWbbWO4gaOwoXshccSPIIXwCf4ODwouh3Gc
M/Wz6t7BNlSgMgeQkciZ00kcZDmQy+A4v1IHibAxkrtNmMYF79sOmhGJs8SPONU0
E+lAYm2ax9ncI4wQC7aRa9BBA1zZctRYW5a8rSlR93h9hvnw4fYqgQXR9bfzUDBj
uUqQ4DE8lqZgsoTrB5P2b7d9mzs4TKM0hK4J089KGsiVy8kSHb2wfN/ugOMSvOGg
wdHmspvKsPFZnjEKIncmg9Ls9Rc+NN5IuKfqT0FLp/epM6+G6lm0YCcTVSPw+Hs1
6Ni4AJteCcUBw6/WnWWp9lwY4/Gcn3PzKixesGUYSPqHX5AnUwftMLAQt8Abpt40
m+oxC4aDb9+2fa33yhbxxmDofvlQeIIEBrqMZPosQc13XALkYEKt0LXnv5Qlkn6v
vno+GCK79UTjHEHsKLSukOEm9Mh5qVSh4mT3fzBaidU=
`protect END_PROTECTED
