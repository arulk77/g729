`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Sfvi0sLTIFcvDesKpgh9GB/PeEldHf9mwTg32vn9TIUm
DcMNQihzXnR0wFKnZORJ766zdUchmPPIxnalAniVuk/7463qjNj3wJAr4RQEpRc+
zzmf3pWUVV5fHjeLhrqRRjGpLA/QvNHSQwfDJRrAjsHx2ROWsXQWe7aaV+5am+uh
bA35jOrg28lVIEnc3VW7p10tZBHpQfQPeEZaHjBigKbMB2h9gH/Fox+6xk2DSSox
2RhG6jTL9YWwZRTuKXQnBv6RqcWSAd0e7IetXJMp7uqgTKH+hD9z61lyfp+tusAt
bIYtqvxkZ2RBFgiA8qiR2gUhLKxdmkmXWoP4OMxxBSVzv4Xx8L6D4uzmhuPmbdsK
xWYpwfAHssoVcayy2UQwZnD4lsYHA9eZeGXi2Ld+n5u+E+V7iWf7EzMFO9zOIEfA
VAlDWjeAK1jwZS1dvbwmO3meW2yk63/GO6hnHgc8YX3ufxF36CE8wjXil8mD3PvR
WVFWsTvDmIAT3qNzQXsxR0gURiab1LWPzJ/TLnrsnT2Ac6owIslZmM2OLTs6tppa
lyzOwtG20UDYmCPuOyOCxgOa4xSmlnw7WGIzs5JHGb2StaDr+7gJxJJDqP0KRpyP
7bsaQhi3ll4oBmVR50/CnRV2h8sfYu+DEyLtkgns6P70S8rAW1n8C+7pkMjOCEAl
BbRlEiIrDgW/SiRK5yhVj/l9j05YwA1cin++kdmCpEOKZPvHydxIL8HcrGIDg/nf
w9L7PNZRus5uVJDBHVBD0Ovsm+tMc7fFLpeTRnyndo2Htsau+bY8suq7SobliyF0
iI9V6FWPL88H6/R88i82H0BGBOpy/CouQ0grmzDBLyvIYbqIKwt6plyV1ajRzhDg
5whkF9SOh0Rjfup6c2SZWg8f7OqcfWIygSkLOddpGLDg+YuUhFAgvW4WNgzsnitf
I4kRsfymnEe8KGDSpHxvciHR3LS646AtsoQu2D5JV1dTY1gUtQ6Vek3s0h5JkSob
56MYiZNVRf6I00Ezv7xRfFrEPj2e9rJWeT0J93HmkWPL0qjWR2CwODzPZ2VKNH9V
lV9MtowmZiO4MEt6ATkpIxVv4BuCIszw2TyI+dDNPjmJcvfwQ+fP0mAupvxvoPKt
E6zL1QrrUjQK3RdbKrHuNlkldFrI0CjypQZ4F8xNZiJLz37/of8WKvYuLhjhbMnw
Gbd6MrrCs2YGLbI9QbsG9uPIoygg+BnaMquseIm4R9uBH1voGbtTnd0JWvyrZAok
sSJdybK8rSH4xFmi9QElWpmCSQzuK0tk0UcprNsnirdTb1Csh4p7m5oj+Fu/H7v3
Xr9KNR2vpxqnmDdz5oD2l7qbWeW1SAUaQbJtOryMo9DgdP4f8AvlhiO+mOL1WnoR
w2O/HTfkBLZ00DYoC1x7664+3fN0XgJzPmgGZlRqOGKO240I2hFibMFCugCRVaIW
zxBLJemtn/t26PLRS2D4+8PJ7Z9qrZeuP5J6g8a08npB1WsNNob6hNDIt6vqHlso
mN2ScPXQ7K2lnujjge7WfpoQNH1Iz+SJcR1Cn/OHchEh6W+PhBevHBcvzPwzcfzW
p6I5oleez6sbXo96bPeL+5D/cm2Q2vJ8SIpdJmxaSqkwZJgNOUVgagnRdA+r8G6M
9reNdCiDs9y74r/PBXAENpXWrRcqgF17SPb2VJyYMtTVraM1w7AjNLwH2lo1LWyr
YGKmOxSEby2c75EQgB5SJ7MYSq5jbaKFXzsO9klx2763msYlD6cmznZZfbrFlaEv
tvMeWkKt4UAjZLEBIL831ykpwxrp7IL3z00qJ8fx1w2lIr4KpJOGeeQunjZBR8FE
bjR2B5COATrNPf1FNGU+z3gfpgJ2gh4jtMWjOW2fyEyt1rsumZM2327JUZEXkUHH
Bb0HlnLm7u5hSoARBtn3hLvyIqou1pyUY5KccpMAUX7xScMMvv9EgteoulIZsvXd
KQVwAzo6Jk7o25onGR2hmrq7SRs5j54uUCMk1fRiISURbDfqGwbepW91VfrsxOBc
VYAfe3I54L9rNORls26oFO+WRiJsd2lbiITvum338Z2aM5KCDhF5SeMYgVTTjxiD
itFIjcquvFRJSTEABtYGn2E1WcC3Si0nZMzspsn9adbcSY8+irTbDAywDNtu/pm9
7hHh0iDO3LIX0gtayc2SOG4oMYji2RLRoFKz9KUXeI34l5PagQfMMiG+8Hq6KSFS
i75Wu76XLJw9GTegVX8Wgwkwtp+sk6EHVxA3w+aPJJAZRftRbdGBeb35EQM5HA7h
4jnYXBqCsktirnpjAUwJzqmoQrfpbnWtYeVT87SDnzCuyseppcmcMX1+cnBMC2GI
tPv+9DHsnQ1phudg89ooze1mC4+m4+TGGNvirWVU0k2v2GxjPt0df+PrJDWJF/lm
Ok966gA3RY+iyyhEou70Naj25vX/sD9mi1Cx8UPcFGuk8kIe+xY3Q0k+Aj6mfG0L
DXujLbJaMFyf0jRB1xH34DHOG6wB0C2am8L1/hQapUi/bTaKFujNhwiNhGvLnmuO
pwW8k1eNteoqWOpufvSLyH/sYD3li2eIxD9k0hseAmBN2iQkn/W2ldbpxpD5BfKl
WeO2L+8eiEhObvEk7KBSKaNz//7XGvR4YL7rWkKZI92qxRjcPRw7eS8XfPA4XydY
8ji54xFS4SOecEzGsvKnIYjNUBy33oGay3NxEWb3xJUBXJO9esd3WdDdX8/Xhi0s
lUmeuR1TQFQmaCNHa249d2oFx8trNCRIW0X8G+IeFFhDHba4XUfckbfu6lcdjXCH
MmaunOFoYt6+1xt6HijbUI1sx0VjCQuLgEX00aw4gPXV0KIUnWeXn1duBQSThweB
CRp1RxGzft01VFkAjky2Uvx01595iJg/FStpwYQZ1e/oxtspxp1O5gv7uobmFgjo
H8u63zn5642Ne/BKe+6k5FkTb4SStEV8o6sUvzXN8i/si9yYr0DcrSt4qxgcqjke
t6WLzjYd0bQstwWnEu+gX/mCHVNNO+sygqBPojBhr4b7sKUNKrnTnhqURTd213Jc
i4aLmw1Wx6LjcGeACy4XSAYxDmzfabM0oxvyHx2dUJxdzOdcQjq1jf9Fyoo5KCQM
cneQBcVtuZS/9bDAOVg16Fze72LlVgx0xGg+gZsmK1MDlo5Ujvwa5lTtSPQnKcNf
JTHtnUq7XyH2f2LRoL628SRrxLrS2LZAiMTXta5fgwrJSvoX1D0zKPcHiMuThLaN
8Ca5C/Oy1n4DEkLv8wXlsHcqMPUaGDNi6wwOSW5lbLczkxnyqNJsjX/QBLOSVDc2
K8sGz1C701uxuLMGL4ZZcfp7sTtWak2zEuhorVuMNUSz5hkkYek1st/LKbEgMIdT
WKdw2KT5ejLLAStgrZ3QNQ==
`protect END_PROTECTED
