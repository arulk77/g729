`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN4YXRffB/CAQZmAXYU593E8lpWXbXxJ4/ZneyZq6lK1E
lmKktXsz1hJTuKDl+MfhmMaGK3A7hfz62qKc9aqmwnX+qug1QSmUDbj977/iL7D/
XnSYY2IJBzvHDENYGmQGkMCA8HuYME7eE6QrhYBZ8d/p/Chdd4ANHbijgDr3W/pE
ia+cpqZq6L4ibGsUSLh3E0Us4CymnL0gwwhHa+7HlEc6/oDSUQUntpgcb4lYe7Ks
esCY3qbyTxDad9dRHzEvLl9RnqE3jHXOinZmJ+/gEL06aFOfB5C0s05e9evwUEbi
5ngDKYSCyRkFlRkrymzl/55bGhQONa+wCj/Vaf6PQq1b6svCNlwDFsUZgp9zPw4y
TTllKElOwG8wplmqjRpqmDN9FDb28vTZ1yyRMykMfqlM+2W9L0GfvFaCotHV3TcD
S15krACjstyJUSAup9yEuKICIdtLj89+O91i0TU4uDKq/X0krP6aCoxCwG7EAuzp
wkDwOe97HRipYIxu4IIul6CUiN9PMcad6tPNVpGZA7ENkdkm9ci+aGNJZusIYqa0
AJ8XimXtCQ0shLZ+WU2MsirQdo7ttFeGzLupyzzaNh5okml4tL7pL5C0773a/O1X
LW35wYOhh2pkRiU7FP+U+9ViyXwFcRggHX9iulygaF8PddTMgOSYZyuY+mBoNr4s
ctCP1duRXsfjXyQTUiYdkCav/O7L/p961vcJqLNB5aSuMdp/V+fjwCtihQo1UBRY
rprehCZWPpP15JR7jh8W2HKRT40iTYyaoBCJ00lzOdPhzepx/nFmRHx9ZrL+StxZ
EbWWg2vuY2iNVKzmUNc3SwDINnraxJDO34PbWRgP7Kzkm7GHAfE8q3MNibQjwdAX
o7bbqfiCzCjVe+D+d9KgUHlgTgwLViuNNqzyaMXFRcoLvku3avQysilLBrrmsNum
rnu3h2dp59Il2UUd3c9Pknu0RnC1zHtNkB4uBKLo1zlqnyIr92g7iFOCgNVEuvxN
9PdF1Lcg6UNEe+cRjjWbYk1f+H5ONXDUPnAbHUT9Und2h3L8svPvF0eTktPLIrC5
5Kzq9obbOQnMnsBG63KUKi16U6QiNlriw+usZZaLsc7YS0yWwfwre4fubfk/aL7F
h8RFHwlIusH3pLsM1r+QiN9g9AHZ9xvkV5jJ/NHZD8DIQrpqz6RhNXKA6d9vXXgV
upIVkaUPjjLB1IT0DGjJicCtiNhum7zKOKZwZxWdg5L+ysNwFXrWWmH/YeF+KYCs
ocgjl18K7zl4sAD6gF1ZP8IhUfPVncI3HgvLt185gd1FpSuvptadD9Jbzd00agJX
b/XjC18kgvulZt2SxQDhTzb14AmnNgmvuapXyKbW4h/ZuZxR9smIOv/wLN0TyZVw
n3F5El/IOCOWUDbMegFv1ipCHLt4q/fC99nzeqeUYFghLXBMt/Mfo9NJpJMQsFE0
26ua0N1DWPGLyP4GubFnn8dFPL0ZZIC0Zd01S19/8vUpUj4EJhR8FLRputsIaJwW
qjtcyupNSWkbOSwoiue+3s8J5/WIqIOMzjSi1AHm/H3Jp6Qr6k0QS5q/FX/ntuNt
hFlZoxnES7SBCrfqfE/9/F6G46COwDN/qJsmyNK8iBgAitWZpAMp4a32PiOiivTK
uGR74cxjPtOpQou/5oMb+oVngXvQlAETY3ciWXrnjAjAF7Xi3I/3CC4HXZxt4LCj
B6F9LJOVUswyPgnglOA1JFMcgzkH7TjN7/t1bq1yUb7In8C+Jv0/zuIDsBIv0rlo
MX2UrYTp7LMwymi3YNtCC1HWsp5duTElzU/vrOGRdx+7NtpWaFzu7w0ipg5IIB2D
JYJZHg2N5zFfk4yfGLZsA3FdLjfiieId+eebNFVAMvIc+BvlsNHTOY2vwmR12Gnb
M7NFSuNuJZiDnGi6lN6UH6UG3/MLZhVvZMiJRHYWHj77k7lGvpEXLJjhRUZfuSwk
tD3m9NZcEKLNfchOQkbA0sGO3OtZTsQT5GASSvmZk88/6ZfE8QbmeMnTlCjJpItq
QuXqvOdz9BERBnEn1Idsowu7dYLi4MENjqDi2CA/+qM0BB95gqh6MX+DfeWZIwJB
YykxbzbudkPKx3E5X74P0iWYwedNLysTjOVZ8AFLNUFF8iAX36S5an4eWJXLb8/U
/sZXOHeZb/S/vcydnMhptRb1FVLA/n3mNv0xPjIpYE/l58U9YwUAa2nF0aVUlcQS
TCU6+WHwn6cbAENx5dVZgHo4PBs+OSE7Ad/B064Y+QLoh48LuBlHwhpPR/MvSnxd
VY7xXQaqPIS5mGoc/Qb10g8dxnBiwNg3jca+TFJwk/GQZ8tMrcSlBouwAbAaUURV
BiqdK0usqxwB2WIQYgC4pg==
`protect END_PROTECTED
