`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/VTvfunN0XBV50A7FfjxGCQm/L6VcWoEhzoztqFbhzpqSPn1MV7y6gCCeyC8Os0p
LC4sTKyRUg2bJ7MkW4iISyIhNuR+sFKaL/iVkuUiuqrmNWerqer0yA5zfv3T9Z1m
snzWwcFdH74h8r56K1OUtgkLkYmaYiVzidKPCs37bCx9GHHQa2Sa39gmGAFDkifN
QYZa9acXyz7TtmU8xf76iLn/fDgTmDFGkqKM5qifJLoi8K7eqpiJWIFX8zcdDwkK
jrvcdRnq+lqi8jpAwpubYwqoU8JkVxjLyRlIxz7Q6b6QKTQjWTmbZHR3wB9PFB3d
tMtclwBV7heGpo/kqF2PUYERXJcqsD5oKQwMdzdIogb73i/8zsOyxm0rCmuSR/4k
2Nt5p99+2zZPH/Wyl0omyqh/XFVKTuydCYNlQoGVMO9aEl4VA7rHW+a+ENzwdei5
SSMT6VfAJ6u5Zn51+s68k04veIgWVkSgdJ/9sshH9S4zi/7y6OttyG12lI5zk2j3
`protect END_PROTECTED
