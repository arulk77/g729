`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIgrWsSZtQVYeGq8+xiy8zsdASlgcTkfenkt8mQZcaJO
XJQFDwFZTqovTVdOJhjzGADIjoQ9L59FtKuboLv2CHX2q4PmZgsRvYLG9z6ZgvLV
k9bX6mEg/gzP6HVIm0E8mjD83pQENiuHYedQ2Owx3O6JTz+DqQcZK8Sl7RgvJZ7w
uzlGPvVI8nnH1QbsadNUcloX+Qm+QKwRqx973CDY2mZU8EvWO5KDG2WulNPHM+xa
or97zNlpRuKlHBV0KMzpQGD5pLga7BvYP19Qs9QxsNXPpvZJ9+1Yc1mcgT/4ntPd
quYB2vPOVOm5V9oNdlB4WRAOxK3gyZNwRnhfrHWu9bi/zatBKiE46QcJBhdzeqDX
ZpQwlySp0Ks9XSMO80hPEgKZBBFfBmu8eSX2jOT7+HnTLsHgn6CnYabMasu3ntfd
lXTyq/CcmfF3dh1IQxgsByystSBig1NC0FsXUujscRIjh2SAjZq0tu2oxKV2Bc/x
yFLmX9bKq5uYWgNoEffD33A6VB43GFgIzIFVDWPzklG6MF2ClroouO21cEM+6PKa
`protect END_PROTECTED
