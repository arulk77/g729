`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu416GZa53CquS+Y3E/0I3sqJvktdPxWl0bGsd8DMx6ZG8
QaUPjUIfFQwgOUA77IlxOYXsitKY8MGwWJwSFAh4XW63eNiN3tQgdB+us8IF7ViI
JKzgOlnA2PI0r6wym/2S/BiveQFYw84jdNKIPPNcMxo=
`protect END_PROTECTED
