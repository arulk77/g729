`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKSu7FWuSXr6W0KuoGvotOANFgkrERlse/eabBK7tFcL
HGFcqB4TmbVq8i9HCuTPpwZhDmKAPaoQzmUfzMelgV4fSLMr6qqnd6iOhw/K2p+y
SieFHUJZP4FeP9J/uG3XUFBIdNJRmiNXB76q6qz9YrmmDZ7kA13t8wdT3207cSxe
wm9Y1t0tWL0SR7CfulFl9w==
`protect END_PROTECTED
