`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4LroAmMWiXymLYBbJ0+dp0mbqqcSWRAlrejPbxWXxR0XDd4yHpxYGBGD0zZEew8V
jFw/7FAYDktLkNOSE+EcNnw52ngOmJlZt7Ays24mvMHSADCQw274837omglgjaU6
9JFK+IhSq+wzADdESuh7IbYLZ9N61+V9xArT51M8iUqr/1Sht14YKWRX758rCJBW
gm/0fJDjncURaOUAQ3sO7W+DYhM5MwySm61GyHvIleVhjOVVoWHTXiFzFf8RwPxy
oCchbvGZ5sddjAjq/ldxSEHS3M7/o3z9Kzpddwgkjh+wHGthpL3uuWNPsRDBnl+E
TbgRARW9xoa1A92GubyxIKATm5nZu3PDpryl4QslHQDyavqjTmbNwMUiJZJGWdco
/cAbcPnBCHXylKUJf8/HFdTkEtkapqKGAU0IBBGJXGke6fkhuHE9oenpahPdHgYE
f1THSU8XQrBNdaYxviXognBW6sHbaQREGioa/1ktjaPE5plYXjghnwq/4EJAqYct
J1yUjdR0OmZuGtQEBjcrlfjmbA+U0dV5nboXseadx51f9UCn/fXxvCqXFTvvdv8u
dEitANRrdbUmk68kd3dibndYlrMEQYoMBkvwYM/FGlg52uXMwdKONg4DzJkEgDDP
kxXLvkYDTSt0OODztWOi8yGuevvaD0cPvwF7B2zMbIRpy5kmmc996d1wTf/w4HGl
mpnyyfnDs46YfFmjt6XXjoHflPNzpY426c5y3unpGiuOoyNEHD9ysy7CSZIeHkNz
jcy8Jzx2MgMUJMUFvEA2bKnpN/RJHXa6UXK4Mt2QsYRaTCPkuAxZLsntiCpLLylL
/qN4UttE1a6vKqv55PyLa/TNHESJK5XFkD/tWJ4vReeUyBp/3B43ilcfjrh0qCbX
ItsUbxQKDoBj4MbD2M5faeZMyeSoa+Gorq1LVIzou4mqcqUhLMeNgJCAmroo3xna
ZjBi/6J+L4uNAJ3ScTAedJB4byqoEVbO6RsBjNvn6L4M7CAmA8xlv0fGN1u5VaV6
gGTr/Dvl93qAEFVTLzLpQfbcDu/c1siykIJR09m6Xt+g7HLPX7ylwjROFUeeZonB
7mAz7+D89m0taihQ2UaYg1bMtgO38RtYeTEEpZA3NSEtjYa+kEBZY31XqXNn1FCW
IDuixWW+GyDiDZv30bYhv+43m+CoLcdq8tFlea0MAEGVGi/Fkvj7dJNRZ2IGaW6D
gnhjuF2J2U8cFp8mLzTI7bCDhMkrzSV8my8E0NePwMO83OiSbjL4OjhYJVZSJx/b
bS1tJ7g0dtW+MCCxNeAU7Q3rvDCEmkmBr3LcRn4s0uRHHz7LFz7/iY99EzpAoMn7
33MpWLnObrcAGS/C0xqYkcnco9QbP7avpULBli/IcH0Flzphee6o0kHG57K2Z7gm
Zvq0t4msIruJ3dkJQF3kfJuqt/XrXGVhR+23FpdRWJ/ABa4wjfNLnfxnplCJ40LR
mOS6qyO7KG9jFsO2Fj9XOIuXfHXhgffBFj9DOQoA72t1Fo4I1bkRcdJesXuBE5Hv
pYltO6VPoFps8CoJKgs9IYLrRg+TMZQayYTZXvqcHN3CTJ114hqoWJ9MA6mjStfO
wogym4xRBP0A08kCB1La1XZSF4ZN6cmqGCmEz+yD0CpgoybEbMBBnazTvQlxzGzj
SlSdMqi8fT+09OhFEMHI2y8tlSmsApZU0InSyqLnzPkaz5FNotojB1kfiYU28sY7
WHIrjnXozJBrpDblzt9BJAR+rZQjoOUOJPNgo5i97LFwo1eMPJC476YCACUdD+qY
ebhJd4GesJQBcUBem6IWDi4Xu5ZbYhSf29HGTA5570tswvhYe+XW/Ra+Cx2QG0yt
P1065hclKszm3HOYe3q9rqnCsFTlveN2K6jLjuVFCO+iXwU2dwxJqtlb00+HnD37
IHJdXj9DLWFhrhddhiHVjo0/tipoDbi1x4BHdZ0nOiRNVWffSkIFAJgfd/X4fFgU
Mx5WVMJpUdDdJlNDNOKErKl35W3RP0SS1yjjQijXDDm08FpyROruWFTljsZb/iPq
RNqs5L0ykfPWhLwTLG/6B4mF5J0O2+VaJMLqw0/bcsnWibcjcF0aLYU8Hf9GjWBc
dYResvIVZmYBbJ+NxWIlPhb4sUBnhZUl7xILrLZlqvN+z5jVbQminvYJtlhKiemn
eslJssd6eWp+WsCz6YuZt3ao6kbGIaWIia605w5UV3yx63hG5rfux+R4bU3rXGtS
ZqK7U1zWKz/ksFaBzfjTqFuSkxjmTi4VVuakuGxywTo+QTGiy43wguIUv2pYo5ML
rVdZmnP9e4LQaD/L1y3IWQ==
`protect END_PROTECTED
