`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLQyxfnW4VF3j9QDCWlYtQpmii1FyPHBuZbwxAUgG6Tsl
ISkdeER39nyNn+dKZskknR5jjff8b07t+TNGNOei5pyeCVlv9qTK+F+mGUam2z8B
HWa91g/nKDTyl2YUnHE7RWrb6FGBkhVSu8/uZYMzORg1nCc+vXhp43QrEkHPKw/c
KZHJLZ7DypanucJnEMAPcX6PX6fTd9a7Vf6qy+wpGA+IPEfSGy7R65mS/12r8aC0
RTr7wNh6Ztry9m+5fEouXLlcdUZNf6z/JpcjADTr9XZmri2K9zEls/SuXpYHOZ/E
98fHsaHoRa50VNwvxsjnaOu3d/u2hkoH+TwpcZlFX8SjB4X/srCgBms3xCJjq7V3
`protect END_PROTECTED
