`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePaUsNaS9DMMclqDGvSPtuqbIog2uyYmBi4CY+JWQTNf
SsU81w4CWaOhmD6rnK2dEvydD4sN8dKGhcTEEykQek/47UYLExJ2NrNfSgp3q8ZB
WIj9wxEVZWfEpmKnUUF8a1zroG/BD5utFmR/iJ8KbPHDU+P+PxnTdXuhEHUM9T77
tP/WU87+YnlnifwfELEmaraLE67mnTlFB9qluACEsjK3YntfHZ8/ZoBfyXwGduPH
WoP/i46NVk+2p58M0TkguhYMeQ7IgWBLOwVAnQ3f6h3MbADAyBHj67P146YNHVAh
sMEicKb8GYCyKIZAqI0sqAyXufIxnNTTgey+rHcUIN5r2PZFzq5f8pJJRfu7+N3r
`protect END_PROTECTED
