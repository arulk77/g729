`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAVExQ+Hs4GcvXmWsTq62ZWB6EqbcspgMIZSWCM7yJ2g
230D0Sb0n279RFqDAHwAm4NY9M/MYQ0uHymiwHOT4WH7hYWt/+ltUGgmLEWkcUAu
Q0O63KtCwR+O+OVKp24hPSqu77360ERRbnAnQKI8+DalwBg+unkcdvErD3GF/ra3
cBCga7xL1epKg0cHOO7rwtRPmXsW/jDK5HKQfrxL5GEfdqNcIdw7pFnRVhANBfhW
BAAn1ZhkVFvsSskW3Qo2jgY3sxXxmOgNx6DV985e4hP2KX5nFcz1nTZqeV9i/jSc
P5+EYX8nZ1/ks2FBejVGE2+AvbWY0J+HunAJ0Qkc5C8Rp8tZB7tED8I/SuzqX1x0
3AtRKxTYhnCNXuZjmA3TlXm4BVxb+SEsDztCAeH6aEFaOTc+HKqw40jNKMAWMzK9
m86Wqfe9jTllssXHK0LySq7TqFUS1NcXw96lIkfoSVkfyMH/nDyIRg020Eu1WZvO
mziwBUR4wd/5ZZW6V9ZVTQXdXpJ7vmk755s9ef/jHWTdw+Qz9FMw3b/R3f8pa22M
yb9KLM5T1BXWdUN0/Cfvp1+1Er5ctBh3DRwJSOFf2Xbe9hAGCznimeq976i9uDNG
iH4v/wFvVQEmfWylx8quToEzbWN+RSsyVqPxl3rgcALhSZxm5qWxbWuzD1nF9qao
uvYx81Jf1ODjSAPMNbX1BQ87/ssErzCtsNKpVRym9jqr075bQRznr0DC5blPOik0
SlVDuhVUdo7Eb362xACeXSxPUE3w6wnczWav8Kb7VJw09OWoRD4k3CDICr5QfIuN
RbmNvGKPiZXJOmC/5f0ia4tTKPzuFTXJ24VFHhjTInc=
`protect END_PROTECTED
