`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB36VS5CZFQB+YDFTuXOGiRG7dZoIjM4CPLSDvbyjZx5
E4wyHHqRPR2PLbJT5UpAaxLUbCPp7ALzr/QPTo8yO7tNE8hc9wYOR94nZ6nMvg6Q
3TTlCCEWvYtKickG6s8jIajq46QwTWzWz2snls4BsTgsd+qIjXuyNI9DeADyml6J
3Wy7jRYZRJ8kiuIQ9jTqG+lB8Tlrdsv1gdDXK1L4fjT9j6SgqB3HS80qBOP2/Cum
L3QbFvCKPpuGtZOgArIkF2AiAxJRqVntRqkeAkw3ot4Y3rdfV49/I9t1fWLQqoO7
/JGw5UX18fl9pzrW71lcmVK+cDcNRf6yBZMYJHRmigTCuY66itZxJCfybPkEgbvm
WNOXVyPKqmu76Eh75EhoOxZoeXHf+GLQJQumJufwZuOY+fOXIHUeDcPXxC+BTP1h
8OuNHp15LG/ekAmr4dM+dZ74C8AXzP+9WDfq11bmh4WmPcfruBhmt2wFbPW9HBX5
7ncLuDkTt4tXgbB5vlx9Wq3JdrbuAnX60DbsY8FJmbcs1R6v/dpEzYPY1FdTQbY3
EiPhnRDnI2uHcgfeqMHjGV7heADOglFe8O+lPwrmQ/mhLyk+xa2tv4dlEKc/n3VH
K0/ba44blDuxz+GT7S8xBAltcOvwySCeG0sxlV8y2Zx0xGUnU8dbvviPmKMTJczs
aSvP6jNqe3am8BlUucSjFOH42nbYXiW9ciIFfooBS7GJNjSJ5E44AdoElIEEzHZO
`protect END_PROTECTED
