`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLR05rcdwupHMtWfh489QpZYCbQG6i9l+rl8wF8SnGaWb
k92tMiH/nepGI8j0rSNqaJ17M+Dlu3AIuw+tLtDhVo/jfvzPnnvbHyF4auKI/hTR
GCpDuLVEt3kZrqlUtioymlgYwF9AZUxAejs/gM1xrLoadtisqLkD3LBu5LaFvWD7
p2Lzj0iwCtQiD3toYq9ziWUb6T0gafBRFKrw78UOrsIR5wA88OQhjEICIntaA3S4
vUEcjdw9s9kEb89aXcu+q+edmPO2S4Rt32EQlnqlDAkYpkYkGQm4vCBuc81QKC7l
jl1+WS7FR3HUDzyY+FV5zj0WJqzRm5ksDYbfOwNwoGdeiHn2SXv8nOkASd8yPq3L
`protect END_PROTECTED
