`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KRHxOfR6PJs4Ird6oKjm1bmyiuGLptx5apfRSlG0P7CVo
tKOTUnz4yUk6N4JHPD5qOg/OnuVvLPVLNQr9HCZFh4LJSLTdvSq8lE4l/gcMbrMk
6yNTZ5eYTnlTt9wNgJ1BiFNQ0/PQzid4otLJ8qIiYnYdL5ZvTQ/UtOkidvhQ0eSw
`protect END_PROTECTED
