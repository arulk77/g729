`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/tycE6sEnfCGAjYjWLGvVX9xSLVIW5qSaB/DaujkDeX
s0OGT8vGdoaZiMEq4JgkX4jv4JBkS9emXBXatsbEjgQZF/FPZ5KAeDwjTI+vij84
fke2K6A1On+6DYCZDGF1XhEaB6vbbdmk9JmPbTkaZ2jlFsop+ntggpkatggFy4OV
YNsLg9he6ETGosapnD2S3NO6Gs4VnQmNYBbUFHBewC12gDdVadeznqI/Bte3js/p
i1yflkk3nnuFalBid02i/ci1pBrNepYrX+UiI4XQW2JKI6YMxNecLFqO69fNldn9
VXdgg2bFXL9hjbGEJXMk9ZaNo+SxnAmRofrzNovQhovpUylduKE0tQdWbQ3yOhVO
7Z1hw1RntJbLUN2rIYoGUw==
`protect END_PROTECTED
