`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43taWTBEYbMBdAwM5Am4UGKj1pMbtHkMCrMO5Kn5+p26
Kzsu9AnqWo3DIMsRZaoTO4thndYpvNYki9tRf4wnSf1tZDBZEcgPvXdviA3gsfWV
khQShQq9NyN4I/qFGZPrleeOGSb7S0cS7KHNpeZveM7djr4QMJV69e5hgXFLY2qC
KRs8wg8k2W9xoF7BYXjNnH6MawgahbMxeVd9HlKVgfOPc7QTDzJFhDdARjj24zuL
b135BpKUw5phmj0ctj/f6GM5rAsY1tAaYcH2VL4HuNm+2RiODYyQxrt6hIQuH+Qd
3wWurVw2vuAgnHuWEiytKj1I1sUFyijYWaHmbrTDIibexjf7spzZwFBICW5/13rL
LG0ATeSSG8evmbhLJnoahQ==
`protect END_PROTECTED
