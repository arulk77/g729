`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48ZmO65ZzJjgZQgKYnDsil8mI0m5O7j7L/Oc+sh756bf
CLZ7fjl6Pwrwi9o39wmyCQbyuxCuiPIygnI5EzPx3c8y/OEMIWzNxjoV+IZvpKkg
z3H/ggZbtcs24FNAo8Kla8spyKQGSgmTGTfaJebXfsSXFgl2o0KfU2+sKz8ItYUq
FwDOS1RH0VQf4BU9OEgBjIQ6kqhYGaBBfd7nLxGrPMg7A/zvR9PJEPe6uk6xYawY
XqkN+/lj2usRbd8Pg9TH08ebuCjHhgWfPVS8Cy7fhmt5LRB+ABNs7+p3r/5IsM7a
A/PTRHExDF2bLgAfNPKyG+tfoHGpvl8FcRaU/NGCTTRDmJW+003qKayJoxNLC1zx
cluPI2mOQzoK2Sg/T9Lj8A==
`protect END_PROTECTED
