`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3cIP9E1nepUubGBK9azHi4w1SUe61eE/ycFSLqD+2xybkRp+SaXgsmiGvf6Wtefw
N+/OWKVqRz2+jAg0e1bQ4yJXryZm3FsG7ooiNdQ0d9zk0tEDfNt9Py3JzARCTGa8
UG9gH2t4HMCnhAO4rOrMsc4ipV3I+WsjHgqeDOCsDTL7R9HvSzd8vyfKpSghNUJn
2ZPZyfLG5BhuqR4XuGb6O8MjnC1yjQT0foD/Aq/iEMTHVO7MKraf2cQLc8JRhb4i
aMSajw48F7qAtNTzOGkBGD8GZ1jh+DYeFs9byPeLxyWxsOYbxnP4ejKbT5/waalw
MEezzjX/kp2j3KiyuMW8dxSrd011YoyAo10Ayg4XedWBncV8NpnaLcx4W6yL3hBL
eGVBajCvhJZpoAZ7m04YBSTnEM5GfIDygh069EAUDNxbaK41+O6Xobdop4J7DIbH
J0jVYI8ZO8T8etYCvVYlaPr2BYfpTiqrMDkS6CG7eHXsJr3IRm4hoiZRS0YIfZEK
tEOugAT+Fz1Ot2vC+3pT2Jm0DTQAaXZQc2LFabC6ec2tO8tnsWVbVwYtPkZjLMgB
S2eUpDIK3SUW2BEfVLbmJmSM5CcilJnHgVOmVY7VS/AefRi+HLP0MTh/HIRj2Km0
49jU9mdzhg5dGWwJ7nOnWkiRebbqUIr55Z5Nc/fcXxnhIFVRtWpYbSUEG727sVce
Cms0biSoCoAc4mYtM2mpUy2m3p4gYXiG5vO8+AqYGl0JqJfp/dc/KVo0gAEO1Fx4
eRJbTECn29qyeuRjOd5XmL0xChZdMbkQrxdwBNf+uhvqgM+nrLPsikSGS3poy5Y2
cnbTGlMeYerHENwu4oeJSvjz+ISaSWXJad1XdXmvq4o4o3gBSvtkFfEMJPW2/QGm
uKC7m4+89vUl8VJYoaCZosPCYMqqz6Iy9dd0QBbnRJu/N7PTPGCvHnFHHOfZ71DG
3/wwbj+dk/C5thxFpUo0yH6J/CnLoVb+K4Wc+zI2+UiHVGtkWeaWH9kTjv9KAZJ/
487XMDANNef+kFRHl1p6sAPwDcxBdEcKFqnuP1VGFXre9ADzZuI6RA1tjTYR3MJX
hUeXwsT7fRGOK4yGKbla3ET/5NzaSSlL/7Hq9ikZ0If/w6Ns9/C64MYrPaZ0ru8H
7izFatoIRJX1o9snuTBzIifjk763FhNqsLMfyjiQjSVf2HRrjDFPm4J1JdupZKnP
lNCOJI1Ec/fC+h+leV9FllPkLlUrI9U0xz+VxTqjR5NMwVE3562HSEX5rdumuJDB
Ic6gWt+rRzTbG1TgYvov0r6o9eLrXiI5VzwEXPkHTbsGgwiu8PgCqBcpztQWytY0
SC5LT/Xzrav6rV7yLkruamlBjbyB3ZzMARqmFPL66b7BCG8juzZzSJswgD5BNiie
gwiwIKlh6u8IwUQ++miNoa+uZBgndTm/4wf9sXITuKMrR8XopnCb3qDNSosDKu8R
X/pGrFHFkCO4tVdQtEWhb1S+cAUOZyHf4nmYNyKKIDy6F4iGs2vbJ6EgzqjnY6gu
FmNuPAq9OuRL//xTfyhc6z8RlKM0ZW6fGP+7VeLfbkhJ5RonjS1VL3pwwgvnShll
NAkVpBwSXV5qbRBRMjLgDELsDChnQVBnTcvsqIvrqZRcWcYY0Z6XuKxsHR5dC7s7
AlyE//QnWXAUTUxdaOK5Btq5bVP3vzjUHzBAdM4i+/YXWgIpBHix2hnZYJPWQoy+
HlvvLxyoTGsxVBAarW0NXXTXdHnDI2ZhWfsSeoDvaxJcmBTVNDjavAiDz07PTrJj
G1PWo14gjPSwLRYVte35humQyC7pyFmcUFMmrpUZdaL2H9MJY/ump2Rj+OizzSKT
kDEZ6nhCC4nAm0obsztnkDEORSYD92bXuV4gsB2dVV2v7YAUOvzPmAwpcFjfZ+Z5
vBHol4DXRG1po9GA7y2LTK8FeBy7xAoz6kX5EtyqkPa9sQIqyAEdJO/ReABw3WPf
6XTzrVppF34Dd8JCwlC/z889iLFkhHgfxJX+x+sCSeH/5mZXq3EN4zesHDJExRYK
WXgWRdDqrC5vpV2/jF+a6MHwNxBUXiaw6z4KGV/L0137F3bjIhG0IIDuUyLsgarD
NZ+sQn7wqroa6YslP0KH0JTBymog85iexvKU57EPzgYVB40n5ywcCNDo87Wl9Xwx
K/Lqa15i8tT8FnOvdvpRdFFRLHhpI7rwTfhg2uK4VWLZ1K8AA7KA0/mLCNHOZGqO
0IEDJdV/HuXQFX8e0pp41Nggb5g330ZYLVxr+wTD8NIXzKfYlg+Sv6gRDDKgJEhW
z4EBOz3s2hNzzVmxxyfV/jyDEaAZWIAP3iTLlGKYnj5u1btJuX/cGSih77P9hy2i
CBYfdGRn78rUtCNZszpezUYX6CJe0Y+pNuKXdmCm14XYj0k7rZDAZwHCFAyN/hkA
yzqng+cUyxdpV+Ws/isJmIO4IvAmuJgKk+T9Xcj7S4HEV2dehykE2nLgmF2md3Av
t4b7STAnCO9R8qy/MvK3wnjYhhJoNdcZPY0ZzUXw1lMRiOElFV592fdOj9vg2TpM
N3PCgC1zwC7ksKHOiLgD3Y80ikZfyIgVo1gtTMagFNQtJEO2zTm2W6zeoKLwAke/
6D9qXPCmrwoVCuZVb97rESwT43puptRkHydXJJWJxgqstqg7h7whdpOugcGweA07
zFNk3PJ32YZ+6BkipSRIAkixoFHZqqwS63lfVfD+7z8ikt84BO+8012NBsTFy6LV
ygYn2Ol2qP7VahnjWrDJN/yzFsaKmDBieUDwhsX8KXilO7okBRvKUsi6l6E6zjoo
e53Xd3wFliCUY8QQaV9xk5lfEhUk9EfPJZVVWRhDXS3FIsZhj/jN2+/VIPzprSTe
jYN4tHGZ9KZiXY1c3A5LQ8pdIGdtb4biulpR/cjMUiJ/H/xFFt8jTG21U0wjTuiz
ng8TzwrD36HZLwCQhH3145goa/K7DiU9EVAMyPeoOuO+gxGb1bli4cOE12hPQLzG
Pw+xRq9G+zyFcsrEAtdee+ZHchfquAMmqIqUIkOnIBV/K0Bnk/wIJaaTdiK1MVOm
Vl0iNKz6XQtBQJHOWoUqSkOo33OgHzSzse/0ekhVjJ0XegCxxYgtcD1oPkqGb/PW
YisDui78MxXDw7KvUoS8CofEwDmFFGpkqJ2AY8dyNCM3zNn8J7WuaccYTESsuEjf
c/3g53GuFlg8CEPcNa5+q2W466sjDxf/wBShVdObgS7jPaQgOjDufqsZ/0NKyFCr
oxn0lPAzDZ/1MCPgH7CGBlBQhd1jDFL7Dpwejan4H9kUWsPrX9msrODhbz0au8mz
41/xzg6zwp02b2kJRA4WXbBBTfJRjAaAlWVmBQEIqQ3rUN731cWj1Rdb86gBhR1r
QeYo9MpxHM378vENuOuXzQ9+48kvnQhYbIb7sHMZ5hKHcRG5xCDPwIP3fkNORZ+v
qDuvQQXGFMyseGf78Y8QfiAOuExc4yNZEDFJTfo6Djf/DGGUNM46XozYg7nQ0alV
wiC0G0caslRR2Nmgqm64HQWMXuMlXZP7DO5toJZhVLf903S11E9ZqKcgDFJZmcQ7
qzox14eU7aP9xgKeBG7etSh0PAL4oNORr8iUDtar2BbLYKd8O6jK/RGMUERL/PNp
JsnlgTWhZC6Qb+aq/EU0q/FsfiYxrl0d2qRtyMMM0mZ7277mREOpFQ7HF52G+uWi
3IONEVSnrkbtOrm221n+jjQHDgYUF6CQRTGgdZfUY+qxUJz8Dm3kxr1VFaqUv0me
08mfdzYRLpe2FaoofZD9xsV1x6vv+zbzCSqKDgMh2xmxer1uQfX1ozrhFoy1PenH
UzOng69WY7p5u6q+ZfveKIRFpQ08sY/rnvpZ9e8jIBlBsgTTTd5SGUSjfdh3zF10
w5WrqYaadqlvFIwTfNqOZ3v2YkrC4r04WFir+EX2JEgg5Q2xCLMKjN3lDGeWOfI1
sgLgp9uIoE9kXgoqsl3F8sRhvGLZ+2HsAci+W/vpV3Izk4lB2aPy9ZN0PXQYcZWW
8ePufD+B6GcKku9NuGCt72lhfGWUh/6AQ4Oyvksb2SBiuFBo9zgN8rjJNTCXbkkx
a2KwZF1+LQtKJ2pvcFVneeOSr5IkAsK9sg2zP7pDX1Mw2ESBlwDvu82HkQ84Fc6f
k7aXFjnhnWmbad5sDPLeMFpphaTGQhH6wTv4GhF9wEvblgoFGOZOpjUEv8Kk2Ee5
JcBM2LXBgahu10neLsJlSutalVsRZRCySF3VX+fWO7olx3Zs7nBYEtHY5goSAyDL
vglXXMrLZhjMgHRVdGGKwzIYrDWin3G+sbJ97x4IKaT1z5FMhVV7kSLoc6f21QoH
KnDQMpWYE3B2pMtVMAlgca3YSMde1RVL5s6g1AZWKTJqBMNMU7w7WS4wcvU4Q5Ot
ZcsTzjC/ov1qN7h8CfBJZ81oWKzofsuPnM8OoNjjdn0f5kgi+lw0Zh4ExrX/fAoH
Xz5CUZqt9CXmVDUivGzs8enuQDf8qJoaAwaDtkoEOb3gyxxu27sUjHXopXPdPU0b
au2GLeNxatY9jog1Mx1klcnfChDJUPj0zgY05jT498+ZLHznJqixTUZ46zgYPfYu
O7sCFmgQ7hivU1l7GzyWlyiRAv9HjnOMj6RisQgj+UFZz2X1szvVkrOxvwPTDF8B
hdSb1CtpEluJYypsfmUMvcg9IEBRigB+2X6kaNzisI+BjIMiyN2OwK4zvKrlF62y
7tMozUF5iqIWob+pSUsueR31cOARoPKdHliit9qhlMaU4/vzH82DSAozEZjkBjPG
NrjrNOuqx01xZGaTIRFN97mTuGNOFePOqGEew6KecjoY/6KBoGOfqo0AQLN2awQf
SPDbs7VP9By5RbBK6t9Mz6QbxTCyWB+KF9FUOgvZ1DhZkBwKmCPlW6JxhH2DyoGY
I2VuIMfvvF3jn+YWVUL9ImKDSbBsf2G3iFb6rZoDI50XYQfKRGTjYd8bMZ64Wx2H
fmRMxtFOy1Q6MwHaT4r1sw4hFDdbuPaagpdCEWqboTaK6WuV3YrQ3d5/UdzqNktU
8Vt6x218AW1xgJhZyUvbcHBSnpyHaq89n81fKGlmJ7wVeYSn9v8n6I/8Iq1Va/9K
0Ia1diKsRQED4njS/Aoi5pq5SPP2A39s7iAD4p/giWtRAzuYH6gSaZWC9f9UCGDX
OdnmwQbR0NF7PoVE3CyLKNAnsX6BMwsRNP1Vs0FImgZqD7sJVEzxq/PGcEt9Ba8F
1PD1oRNpKwHJjZu9wHvmhwuyBobeS71IPc/39ErL4hv0YoH1Y5LNC8LwzDAogtdF
j74CRN9U81V6Hw0OEV+hi5KCMnWJ12LcnNWrd7f9jkvf0jvr4sqKYPx6EUTEknII
VIWm2RvB6fDmc4CTFn1O5WQci1lILPrimIM6WXU2L43MEsLPfWOWIWVOuUza9TBx
y2BEfsgzvhFTBluIfHtNKnAXFHDNaH/xCT1lbhoPWGLywZQw7c4NCT78qS2M2DdT
Olz4JodEP9eEqibWejGD79iuMB2qF4IBNOt90hyO2RqvfqM/KfWn3vOBpq2iJHjC
k5nWQ9vyWtfr8NB755Kg/9QY9GTV8BtQDyykAmG0Ehi/R7K/MO3+4kfyJr0Jx5G8
OxCoJ0t4JHcNKYfvW5B1lhOU/CAyc6TpSOBipTTHcTH37qoPYIC78anhxWMSj/zy
jYKio7qn8K9pMCbpYesDjOAucxSfpr5gxq+g3sEgpFqksi74ju+BEzL61aVgBa8e
9vgsfstYa0krhBiTdsxm+HDD24Ma1buVijCUoi/BVnswxTMe2EmlhbpA7t8yrH/A
b2dEVVZoSwrLiahnywRNQuKaJXJ0Hgz+dBr99OtZAHzZFmabggfoehICLPN4KrWW
pCtpbCnDbIfVwqLqF86YG0/kFzNFMarXabFeurqxY56P0gaHkK1Y7M8ltZPX413r
IUkMDPu2yG6A76FvOygCC6/9BCrbqNYLP6HKb97EFJk/scEVtRL872dX5BG05SpL
uSLf5F7hg2rm/GxINzXiXZPZkUJwvkXGynk3WJPtAF3pEsEXfkEhJYYf43EKzcg+
vyhklbm2sQARIPrjO3TRjwROX5IDsmtYDWXL+BiLCQvx3p0FzM1LPEeWkPuiJq4u
NYXM4iNsgZqeT1wC/ziOENFgMtB2N88ZsjLKxKSWTj8i8vjGpacU5rR/VZSxl7Za
IbLOO4l04qlOQEWsXlzx4l0sf8JO0zHtHwFOuEvcfhMJY6xBkX4uSYs3SDYbrFEg
KOxhg100o6krYd3Al0zJDYxec2cPYsPkqHjt2uKpIfdQBPETeVE8CqFDrnUzRTlk
9LrOMO6iUwEcURII++P6VQbbWyfWnxe9k8TtPIydfKIHkQ++IyNgbaGc02o/6HEi
gQe1DMwH8fBYu64h3CcIH7oDUcOyyT/EU8AwCEhJhlfzPaIKwnToXxGJhyw5jSB7
IZU5V8g5eTnIclcXFFW7eRZ4ubF7og87AuSgxzNMr3HInVfGdLJm04xxaCgWJbfw
9pSqo7MZ3Ibpg1LYPWiXxThJKutfoiaspMscXeg1tv8pZFwstgn03xQcOiJDch/5
Bq3Ra3E4k6rPqy+2l1WIA5u+FAr4HprQuxl+CGXIpKRYypz21EPAlTGZH2fP3U+G
QB20OM7u36D1Hy3kRPrBy/8LwNrRrN7U6SHH4CzUHOhwG6x9+9SPlQgOzw7Qgx1z
JnVyRsC+WcEt1Y62cFQx4+FiaSzqWOoobQbcGTb0jDG5L1jutxhD9HWjzfaE/laV
2kBEdMunSaLBdPjIfaoQalbMmOY/0zUyoCxIFxtqDH1nDCSzlFnKUTlvbhq0IdFe
gyQjYCsJjU/lRcSN1V35mUsN7cYH4FGIQ0Dxd+CaXkJk+7aBp5xHumuYYrUb5ifj
dLtt43CMGxC5XuC/WfcWb+OgHJtmHb4TsyM/Z8B3sRK4fuMARW6KxMZqOgkGgO8O
QfiFhENFhk0N3qjXpe5/KXe7Qn2G/kHHG8RvigbWjX79mY6Pb1wvSCL3bGfmio78
vJQxI0L0vw7lEuNYzSIX4XqqY2buNzf13U7puHP8+sqsg6w8SsXUNOAaxeI5g+LK
W53S4xhl86hJM4vipUZyerNkPG6iIpSfoky5yG6t4zQrOZXleI3fx9sDZRFSwpIU
EZHVwZFS6iHwlNEYEBElAYLeWS18cKkV9DddugoUpki732DFoNdYgns6cLu/L3cA
QMyHcnlXUYvl/28DKJT3vnvjsFMY0pNKj+qGp8RsFE0IWPOydluzIIFgXPjTp2C/
mLV03ruJhqd2u70xR1yXsLdaQHLLoy4iwvh1HBykq7W+T5w3w08m1plxapfnZgi7
1+AbZ+5FPBwVF4gLxB1/+/pm0QsnkTCNe+gFgZcARrQbpbWMzlz3pqsTXJlLgCOJ
A9kkNtrR58gcV5Z4Y9axuA+tm4iM8pc2GHYhTEpsoT2fuQUanVp5jdMUjxqb/68v
5xR3tiKjlc1G02MMimjzrIDAsHCGeyQ4zZReonIs+AEYKRfTpTr/cdFDRnpY8JOg
ZudtqLm8TkbKdqH7wUmfuZVXXecb+iksrqHlTxDDC/iHzG6MzzxY/uTFw95PkVIp
g0Yv6g31Vl4w5ZSwgPcjVpkRt3tsnhf0mL4Wl/L8SGC7xRHa7hErt1UvGKZyOiP0
3aGl5fIJmnAqeEcVCbQljPzBiZN2GXgdWLcRe/kGSpMmsQAEJP8/kYjOBf66r7rS
n3hdWx0fVpjCAQtf6HC6485MpyiZZbAZ2A32YS71i/17CYJ9IIGieJydnUk3EDRA
5o04Y6/MSYppt02Mp4rcWqJld3V992PLlnY9YMaZwZdS/941w+8j6TCaY86w7Pxw
47J4hUVTgjLqM7XTLbVrATmMIsZgNNd1uhBh5l090eVjsvblQ7Oo8P/SA8p0V0Mt
Rnci1qRSz2u7e9Ij4szffIKg/R9GzfKCEk+iUxEXftDcZQ1w/ePbB75cnAaWMjaL
5YOCIfgUVIUDHeQLHs//G+x3BpYhuD1HuA+A4NJWAo5sKxwF0GesejpOdX70iGh0
mgQt1tbAOI+6coT7jYdKT+ii1YJuvRH3SqXdFBiuDFvdLxq7B+B/leM4zGMyZWU+
ebLhWoj/glzEyC2MSGR2/MM5EmY0BWHSvdPUXRUGgO5JY1N/ReKErwRk3lfVW0pc
uFbD64ZBHYGC4HqqiH/9qe5iaeiFqH0NW1bEFCTpbw6hQD/bAWqonYKZG4loF9fT
YFrIvLiPsoRbAyYKwrvQx2MlgBOlCLoVPNdPyVpUpEYuZJrutEUNj2MW0N6/kZWF
YwmdsJXgADXhoteOc+1BzexkvGuA/H2d14BnAM/R3HZXqYjTIBgyZpsYw8q2Zu1a
VGXugbmXhaZIC2ygQDFS6btK6OQAwPllf/Vu0laZcSNozF/ePg9Ih+ValVKK811t
z5E8UjJAs/cMGCZULKbMDwdTIj/FcTohYP49/k2I+niITelcGuB916YWWHSVDqn3
0XHJGS0T5gz2+nq9OO5NnEI4l/fMmP7SPxGVBkirh7KkoLmGpIOFHxN4eeweA6wJ
1YW62nmbqSAc6nOjDnlJXL5zvi7uGjyGNDXRLXcIjmfuPQbzGH5C666R2EqPhqjy
t9ftTq/whdDbeTb5JfFzMaHLq3yK2SEWIps+B1IYhT/czY9MjokrhhVYe0iVQNTF
t2sOQvpeyxPtEdJaB2thXdySZs6QIf2VY/PQtgXZsWgjHaWCPvfJFfe8u3tDyD8z
u8em7fj2zL/Xrb1T4Rbzf+LThHsw7V0fiA1M+yT8/406JLT11yS7oNh7VgcMAo63
q1+K/nuOn4T57Z4ryZFgifWEDtT0itdGWYQV03a1Av9U2M/cn85lS+yVc2ZI3n3+
JADAXeVlkumSxP0aXsEv0mIc6+GJPcMzb/rkCPYawy16Zc8erU1x1WSCVYCXoeWK
dWPAIZ0/M1o8+KAP25TCR7cttTKhfp++qe40Fd1ut7QneclAscd/rgt7oSOfLvkU
uAmoKdAjsn88JVeLIHokKZ1Nhv5qEe1QDL9c9qnSCmnqFkx52yqD5cnf67xRQ9PM
uzE50Iv+AAerzrmGvGV/lLqFDn797R/Cbw/GqqpundBYq7pXPk1s/d82/8F0Kk2f
bMFC8aDBnYYiO8oUiZx2L5bdPQf1lXiW2FVyAAg6yBnCd8xho9U1QQipQ4fFGLph
TRzyj8EtqHByniJxC9aKwfczJXw+htsWeS30d8XvBOGsShSnyYOgpNkDYzu47x+6
odo0ffqf+E5lQiOTg50oMmnQeaVhtINNZ3/AJwOqBn4LLNirngT44toCYzuFKwk1
dgfsi3BdhBawqNAqU2aaMK9ip+EE8mvQ4w988GddDbzpOtuZeXdB9wRDL7dqPGok
2AUW8penDXaVYUhvN6WoU5mlwUeg+n1rrv8Y0f13x+eozFGZYH1q138ycZ3ZCUJY
yZR06TlnFJSI9hYxVSz8jzgFRWXJsFiQCPUUW7p/wGeFkQ2EDEZj/P2+OlJyU3XR
KqQaLXirolzZrTguJfcQeTp4rzgof1Oshd3l9OevK2ggPQGBlzuc4RkHl5uSiV42
nH8Sn6fm9PggnDtfnIQVPWrenLFA6xmEae+O0RQDdCjWZKbEJBc8+RhJoOpV3Qb0
LFbs9mzCNW4yAbo2gHkL92yGHXdjYUQgE6TcLDtqGCPwy5GMdLc1c0zMfoMzF+8i
WCPkt7RrUpw5vN28zCwt6QtNZnBgWsBj9gNKB06q/xiM33XjDuREyBenrpu7EuMU
81fTM8Jmrg54LXva4joSKdR0eaEDTg8P0JSd5KvQhiTTzIyNgUqKozMgn1ZiM1ih
r5W+uxJBdwlRUj7o5ACXYKKVdY70/IZqdVCw6rWLOZNY9tSiwU1pZmuKNnWFRQk9
+5ITGwA8ZTaORgWWIIXKSqHhjyFoGZzAef3eA14Q2RiiNiIw2PeJwYNsmqQJ3+4O
ep67IbaHJkTqCXBnKK21ul72PGW4fZm8CnOrSB5dfR5JiWXfQPGsruGYeBMHXb+k
QL0XwWIiZn8OFdlce1lATKhcOrYi7QsUCmpUD2z8JT7Zt0ZiN5yJIxWV0pbhkw3E
C/DKNRLaWGAqz0nnQYSN4oNCNy9gD1u8+ZFyqKBZeR2VgIB1spPU6brI80CzuHIJ
CL5HXpfePZg5kpepDUGXC26nf28foNr//9d1PD0MR6AOYuzBpcggr1qXdTfkm9Yk
t4KLQQ7txbxswyfsjJfbh83oXyIqXjb1pKOLgju3+/N2kspo+Z3Et1+46Yx79OEU
D4LIv87a0ahBAU1QMMjsxU0+Wa4aVFo/Yyj5GCDBc5gH5LIt0WI/zgAyUHGbWLAM
DWJgu04vEvwVPvC4vcb5tf7osvKb4Tcg93FAhy04tKUhXH0a1rDmsMiU2tnzUJ/G
F5XlPFt+HxcIkVzwdgPP8pnpr247Jw0Ya85OIWWN1VN7DhFzLZ6PSFcTrEQuenwf
PGx2RbQyNPInBslwI5fDoxXwCLeNd2Vu16Td0bLLiZmh+OGjRuHPsQXHWvQWqE7I
DB90u8JGW7NxCc3hiqNVpfs9kqTYsO5D0Xqvr+3wiXLXqETuB1WBqPTR9Ztct4e0
bCamjRabmu1fKAe/C13NmGJd3Xwdwacb9Zyo1CGLl7vXjD+V2GnnmBJkDkZvjxkZ
VqgBMi+OXhtfLuHkfJsmFgOmlJLlC6qUMgQbJV+R73SIQmbrTMt8JfHSc7+TAKrX
0Z9MudBUeW1AV/PfMt72tCATC10bLDRf+aRBfV1jqKn3c+RAz3zJxe2j23J6Iv/n
qQ6EMtKnguh+k+3L8ZDxH3WXnFLn6djaFtwgOWBPe7K9in/pUzTyNHlRWSogrqwb
EA2q7uY2dc5zeXcek9NlnHz/YDvxANg3CodMdAg9WyWC13G0RKkwQVo3hFXztNav
z0jfN1jWp7ycblHjHOmoyzNbfLfyAInffM/2+Kl7bDcmEHdglD+kl34ELHG9KZ/S
VCIc+KKuQkABx3QCu/IfL+KKEhL+KfiaoAFgfjDs2gLE0eAI9zhZgHGKVt1+MFx7
TxFJ3x0d3DmD/S/YX+kZ5chgmpq6pyeUCsgsvlTNHtJSAkKaLVzCsWZdfUVw6JbF
3TxC8gjPwzkCAndAzOn6amp8DNTG7wu0HnZ4dltUubYCHBxQ3b+S6OadGNWXUd7R
/4k2LkiRLzUjmkBx28xqFjDMBF18ly9izxNDNNeeACL2jgjvx9CcE2i9dh2yYBXh
rxFvOGbJlseQ2iQOQ9qlADlwn89fIzfECOgex3kfjZjb+GaC9CbB+5ldOhwbMCJQ
Ryyk49tGq4VkcTiEdHbfpECcHBYcCE3UpM58erWvyE53DIzt4M4mrmlp0FntJSn5
m1WqHGUMH0GaD2qKolr1tAz9barnX+ftUjKb/SM8/qCW3w/saH3PorVCjHIiQb95
cuXr5UaAPRKJ6zOFjxLQad4G8GA0daMTQrtV/FActuSzgcpB3YhEMXiokD9rCKul
mKhxysMGN1HRLHNy1lByH6j460nN54sIQTeXXrgIOmE8s/Om8Bfz8vG5DC9UVWY/
ODv/9ZoXUbxIlt98R5c9Q2jSRUJhgNYV2RsgDfESsI/gzqIjIH7vFCrUDMhCxwjE
q5hgKuXrZdz9XdAxOtmwZ9SKDnHphCSWnA9genW4W80QbkAksVohfGA2wfBpl+3v
O03jQCZ8pN/ptuy+R/jzwcta3zkOvPhufBs7SiKN9yqrIrWO+lPJ9cOYl6OQ1lCJ
edFYUIrcXJ4iZ916SXKPbZ8GX+2HJctQnmR5OrkcTylVa2io+4oLT/0Zqby2+9fN
7+SuAjAL3W5EmiswAeyxryG8yBbxGG2YNomqaEd4WD8heVL8c3HKgl1rUsN1JaGi
SqH9TtUWlvBSPfpEekLO6FRm00I1FYA1zhn5D2YkL0Ok/RZsjx32L/s24sTyoCWk
zPwDWAWgNh+EqEzWcBlS7Eojfn/vXcBXAasBGdJE6o1y+lDEuEefezOEOCY/CeIc
Gq+DadOwItvv2LoS0T/X3XxsX9hPgQ1emPYvyyoBb6BW82L2b2fS65mw1L8ak3rl
7PSbFxIozMuM6ueIwedTkRWU/E+FMvs94OaHGepUIcCSLCLdqQhQgB8jzVY0XhgT
heRMgsuhUkaznsNZf+DaKMsx5R8UZMcXWyO1GRc3Yazc+ybUbmlK0YgGikO2eEHr
G/dE+KwmTKXxmmybCdzgQPArS5ADEYbCA9egJx3v4Zaa9iytK9PFYl+6+3MrixOR
urtJq0sjC/cnrNVYjOYdaYqwt6m/+O2sfjwmCyyaB/soel55UDsREszUFfdFTCte
cWkY0m24CwZ8oVJYFGF6uE+mG8Iqkh+ai3/OqDKlD3Mwg6KWZQsfIF244GZwjTi3
xp0OYFdq08FAxpXuCO6MSycrKj96N6/qiQc/Va+K8ngZyB7HLFzXU+MNJElgoWFx
39j+I9awL2LVeZLk7Qimns942fNsst3rnigE3AgKPlqmc+lWbeZab2JHCFxBOBRC
Nntc4l7ZwPGDwXKREzF98jPHn/lSQGFvL27AHdlydhGk0nwjUV2zBJP9/iSE3WRW
znM9sB21goepKItr8hE7Vca5bgWfX9vkAJspoWXdEx6YclxzO77IBIW9BjVDNxk3
`protect END_PROTECTED
