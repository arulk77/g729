`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rSLajklFVC0O+X23/xjtlTaJEEpVFvJln10u1eE8sxhFSrKWXsqWqBHzpoM9vsCi
yhOkf0vJbAmRt4OxMC3fW1U8/7DXRUQr7ZeAvnp1gBObkijMd3506L0Ahdam8DL8
0+5xlIYCOdPCJujLH3TIpb9jpST7K7af9bhbGtJkm0u+HqHi6WhMoGT5b0IcMN0t
gtE3wPFHjeyp++GyXlWnnfPxjr1f2ziKY6Z75wLdr4px4saCHT5gXRRBvTF534s+
sNsbidaL9x6Bpc+zLRbA3iQJr4f+WHnMdQluRlgYTfs=
`protect END_PROTECTED
