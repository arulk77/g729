`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zduGlkiGswLfE3JRjCFQ0IG+sGDb+yPTM5tpoEj/LRt
nIZzKvRc4BO1WwB55HQeGDPzxBduic5yLNUhe2fBHnaGb5I1z9Gun1SWJoRDqejW
ms5ramUoMLVgKgYlICnHArkyDaPwsqxw1e5SlEtRrTM94TVgXyX2hPMCwyZLNVuM
vz3TQ4mo23mgiL2FlF/WmIGO8FZ+EjL9g+T4kMMtm604drD/fGWQgorUW849TZiW
ODX0EdZSZgM52XW9FfG6RIv441bc96tqBEfCge7IjjR5nebP60GQ3PgzpM/HMG8J
S12WIYtjZL7DjOtrtvn+VA==
`protect END_PROTECTED
