`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHLohqqQ5DNzlwoh2lMCzzbwok7Xb2J07V6vlC8Xtt3Q
DdzK6m+UlB5tvjToXYI02slSrAOTU6+mUMRQtDEUhD5MQ0IIAYzrDXKbOzwwvCI9
M4MoqY52MVWvcvmHuOY3sx0A/9N8824OTNmwDyuSsEdfov8Xkxq43S29NsQP6oTQ
1W5CeNeFSGHkDFEtZ5/usg==
`protect END_PROTECTED
