`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN+E7q7m7XNb48gEKAyCOpeBAdeRhpv4GZsAnw3OPHMgu
mH+r/H0AA+aZXwMdzSityRpkcHjhajE0IrrOBs6lFO69eHuTBjkDln5EqOZEjA57
964ic1BeObVZ4pLzQGfLwoHwpmdv5dZ49B8kZI5JIiBbqO1lqbFn7m2+wnZUrZzB
a4itQRGNTTMrfub+pnCA1gUSv/h/S8f8XUZB9+sORmEcrlbfXQzVex3rKYCB5YKp
iXrQMt89KuWHWI83Ognxccwk3o72pjo15YLBOSspIsmvoRFBNLwsawZL/J7MpSyS
z7t1hRxXXoaI6IH5ZBBvMDmEILFpqtD2Wb4A/6zCOtZXI2YkEqsH9/FU7rMpUUqg
120dLBe3mdg+/DL7nePrgFiN7iN7dxl6HYux5kD+eJLPGbUYlEOMgy+xtzgcs+1H
goLcEJObEBIeO15QI7Ch+2pQOQ133k3AiJY0fom3HPUTjZ5wHfbwG/wuDyJ0IzPQ
xoroSD+2HEr8cZ4LGXqKmCph9Hb05TMLF7kgNu+3+JPIpMnaNV3Ojjlv3SeCPjbD
nqyckFaw5wrHF4V6uV5txl6R7GbAbdzH5rP1xyWUsg5PimkNMYVt7+0sQwurtsvv
gC/kodqraVgEuhuxg96E93oEtRnhiOLredYiGBwPolYZ9BWjd6+SMlPUTIi4s4BR
MHp3UuEVxp1ZXrCZyHRtH8dUexxryLGKqlT7/VeEDbwwvN29opd+VvReLKxdpDTy
H0kY8yOrEf04FXxWOwQQqJnbyQrYGfE1w7GlS9617UmMRDdFJgkkMiihJqczsKbm
3yMBiLBv3kKOr0wK4BBkQpTdRLAyt0y7nt5eMFfjSgvCsp5xM+rRZ/KMMvU5RKPf
JhWwtrbvrUBlB8c7nAZa0w8qA3F25zEpCk5tRd3UZIpvpC1aOqo3jWui+5f/B/XU
sIa/0DKRASg1MmUCo8Esd4ayQf+H6RzjZp33lRmFVScgcRkHyU6z+lG/nb5lBmv4
TbyD6Eu3DN23tgWcPLjIYsLNdjiXaRziTKdqMuCC4AhTvcyahHzQszGEibHslUGP
7924eaXeKiCit6cPmQEARmkoODMzLlZdLIfHDZkGhyKVYRZ1AcDMU3CWJak3EU4r
yGP0UPcDOfzCiNi23wZzagdSNhqZaXk7/GWkQxOFDZ89uIQjSGI17uZK8iJe+5Qn
BHLTR7cCVuHtCY3b87vh1gEw+ydiZiElP9yVQo2vWlwo9QdedjUj03Tpvo+6HhOK
yboPurSLZE6RDUZvrNfp0kN4ZKS2KUHSLUt613SPIF1DXIB4zNaTBsq4sCx0YS+4
bmwr10gMc4t7d8ISBeWP4g==
`protect END_PROTECTED
