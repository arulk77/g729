`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SSGVEcuEHKvxmSL0nCGALMhx2wUCSoQZmZHyIdZrmmWI
1/DdksZa2bbKxJT0R7t3ha2+D/jfMitQ+WCKC3KHNzNIHBg25b0/vSCrJVKh+tFC
IQ85Xk2Kr32Gtiw1voyFXh6C4Gf20tZW2vWDOzZ331E+rIeabIxOpv5xiYUC6Kcs
LNcpssCINBFxpQBoSS2oGwhTvrpfotSI/yyNGX1RFLf5M2x0TnupY86jdizQowZX
US/MC+6fkUEVozTUDhUb9nG/0GHruS4OFzphuwEcucQXe6LJSTiStEtiBWzEn6oy
8mLd/tVb0ewm7sN7glcQrRukxUKipmVWQT8Kq0gmPOVeLSH59Qo3BjAhij6loZqg
bsNRWiYzXr6aPn7EuV0uWekWubgfEkp+NJgN6JIuzziFUGCthKQS04nipfcRHk2c
/CRWNR53RC+S2RBL8Pb+MCseQS4fCpw7mN6sEpgAPjAhsE8OfTGc5enw+V0hDXPL
UYpoUB1RUZXea7slgBibTClYJ6uwI1R4LrjwheTfR07vDqdxd+fA2xhtsK7NPxLi
OG6buRfseV3VkhWLB6RdX4sfX+Tl2VluMaRhoz+/abEAh0kG1GrBtCJLOodlDlMB
x7nSAU7jt7zX6KBKwXds2qdyrIzpVPW8DAX82uKMqH5JJbmfEI7sMzkts1Rgxr//
Y+yqwTjZDL4OHXjYdxE2TZHdGIRQl+CfGrbmCmoFMK6p/MgpdYkhtDqHuK3k4cul
zhlNQlrhyB9OWy3INcVQ/PHeNTaEa8I/M25nDW2MF4fjIFtu2f73+SJQR3Y+ARkW
7l/ZGUhsJIrXFlfAEeCAig/Li5o2QZI/XFhoiQBKJiVatHnClnbx9okgVWML5uHt
Pi04lV1ItyAam/tfW4VgIonoDftzTWO8oOjJUSS1F/OnPuBxw7Qev+6v+0B+6elY
aG59HospO9ejPlOnernRZMDwA79MEu6lzaUIvIzDAarWH/puj/r2hd90PY8tJm71
j/8w+dnQAYa0hq3HpXwtrs8hIdujQDxRw9P5XkVoZOUAdp0aEpMGxBSHBcS3KK3+
+k42GI2RsxOJimRhrg0QJDiXqiP3i2dvBQ5lp9FJoiUErpEmerdGtKYp4lkS7ByB
nTvcs74GL+bU48ymVIoqmrAdAOr1wYHzNP6sYnx8x6oWq70ahh1hLOy+PbUeUW6m
dYYVr1A71NjRygly4eRgIT5kbZT6coJeRhxx+tzgokp/R6fiWP3nrGYs79212Qql
v/e38F20GBWf/3+1uDB2gJkN7635rgTxe5MZYoxo1Bwa6w15IOC5X4aTIPbtcCyl
1Pj7AkRAe8Ln5jySnpuZzXYWUHjhkeriwK67ynvzVrcXtu6AcxRvURFsSu+Go7tF
CzxztjasksdIVgLqQTWYmqhw4hYAIJmLxu0S1XXUh7tzvNgjuSxjBckl+JWRS/BN
NWDbAoEhsq/eWBiAlUZU66mhM0JYolia84kBTxndI6B1NAeWjREswHSs584x/kPa
L/kPXKEwfxbMpabeqwHU5fVRWEXdSLl6OzV/G9Ob97LO4Cl5sOhrkMZvrHobKnM6
wGsTCQzIUce06z+KNt/JjBKnGUTkFLrV75KaKZKzaXcYHmdS/1D9usfkSoakZOrk
Vo8Z1uIdTMZzeofIf19j3w9zS3SKPn1P5eMUIRJArMac8YzQPhTP4XsGxbhYfL/h
DzU0iG5SO/7gWT1vgmTNVvRQwUKzT39zTOFz3UgcRAyvzpC38fv4WGFBbbTJ72b3
qasgk+R67TjnGekiXr32TCkb6X1v6Lzeyi64DfUahGHHrZDpTiLkMhguQrXTYfWh
8fPJsv13I2pUWWW4zajZjLXZ17UgAGnN3Sr3Ce1HofKXOR2J9cLIN87JUb2jw6K7
rpyV2EuyaVimBqxo+qJAtIbG1K+LfRwFEZwTuuJG9eljrBQ78gmzGhxu+1kI7iNe
SbZf2WVHYHn/5PgiJS8+An/yr8L90W87BtI8h6tixgDege9ujFDcbiF36Vk0Mr/k
wJFpZ4HMC5O7x6mZygDOWjeRkx/0bjjwTP8o6pcTAwn9RXABMSHABNMD+1c7kEmy
4BuhYYzmUXYDAYRJFpYZw4YN/YIrNWKuX3j/zNmzGK9yBklp1DoStoh7nQQjAiIM
Ocqgs1hJ4hcw1XNdS/bwQYElmC+CnN5RJUaPI7q2STrIpG3NZkGavY/tQwkAtfIM
l8rzMHLB1u0/gTWplf4SWJ5n8UAxNz3H6wMudFn0EAv9iZPSwyFm71V1hrz9A6I2
P8Hjzfe8NbniY3Vd+Ksvgamfq7vBeV3bUYEQP7w9iDjeq3o83NjHB0sW/9TzxMcP
8/DVue4d2ako4g7Dj2hv3uwZ8quT5l1oJkCuZQ3hhcaGJuebwVK0NK4GPpqSWK+1
I+xV+hEoXN4Gl2J72+tm5l5+n9JJFDqQe8o0tg8wc9A1+4l+G4vq1MlzHEXl20BV
t7dypSQDV5WS7SbjHpEVdknJbT9tSIno7EyIq72WQO6fMytFyYsgvoNg4ErFxcDE
BW4/BdTzEjAbmOqLGbsmCurgJ7dsckPnu1lzJuzwhaHeYaB7uxJEG+WO8jR4buk3
wgv9uJ/lCTeezNF0pmbEq33jAGylOjT/IIvd+x40dZJZE6HWQLlp3qJcamrFFGeB
1t2wcyb+kr/NnzlNHu8a25GKmmBI6M4QfKftucrGuC7DLiKOAp8ZkM7oVXkG8Wc/
qJa43Icg3qKR2M1WbZYu38IzoXqPYTEvlyfe2+DPzH94JJqbPwqwN7ijLmkXJvH6
//JpJcJXut1bGftphAHU4WiRQ2CWrW/AvbZepoYZnojIybptR4zWI8rv0dCGg2Gb
wITCPl2mM5CmmhKCaZmg7poMzUl+H9DPW0x9LcRSv0El3xk99Ipdmcsup0snoUpB
rhE6yhB1RHWKuki/rcBCCYSKZ20UDt2+9qW354nnFz0KuVm7Udoi20zbhRgVK+UF
y3p7chnkaVbFW7bEMBDPhMsK5AaXKjTd8Sg67LtXcJ5yZ7mY0lkGXW/FEj2qJH0m
kLi5YwZSYOz/iqiFe89p5QOo+vr48BLEY/yWDD6KPZHXDprrRAT3zl2v7NzLsTFU
R5+LAjqNnqHlhmyK8eEWd8O6LkOvrpK9DbFXGcYPFD79leh0B8n7Zb3Z7VUjsrlK
y4sx5C6Bt5mF3PQMFarL9gJMcCL6UeeXOF94XG0PeSvYum6HuW/05hOmyv/zo6Wr
Ksn0VitZfeytbCXWBZn1Yg1hKcQDmQDWRYlnlZusmARwuxoeZzzYjNhThYWYpDgv
XTGpICHhmYQCEwh9eiHjmYIKS4L+JOpf1XCWOv33Fqm6DczzangXxxQBBQ7zvqXZ
9RbVUq7Jh9kQF2Plr0s9+6W3a274eMgBGs7yiQGwIDxY4LVTEMp4CGTx17MJBtE7
nNMNCzEYC6tida77oWEM622CCmw7KMcd4VGLlRMhTAPq+aulkVdMMsD/E7di6Ihm
Fx06xvpUeiKbKyOw5dJfrsBnjCjR8BnMBSd66lcbFdQ3N+3E6YmWcqpHU0wbm0lC
VMzDhTxNQSHfVfqZO0zmmuv+eA3enCicPxnLd0TXl6w=
`protect END_PROTECTED
