`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFMCG3FUIxOHGkzhpYGfyBpd9vZR1LIOFGovvr91mX8/
80Cb+Df+UK9SUteIUz0YrklGPfc967QCRX3pBAk5yH0EerENzF/eYgApH+Hy3Afl
wCi5AHY1EPL54xTCwrZhOlwvt2DLuERbb9XDuG/5BAwUEDY9I27IhoscsEWYpffa
MUBYFQS9CFd30QhT4xEom9/zCD+PKvUD5RkKujyLGT7KgkeFrV7RF2titjJknHtL
opt05AiKJiiMHFcy2B7N4VvRMmcx3FRi1mwseNow54l+Sk/vtC/DpcyDtAQFWKB7
XZCwrvPVcUT93AW+QPs5ADsmp8nb4JNeyu7QlJTqjWS56C2mN2yWhZ98+/tg9pzu
vr5jQ6r20qpWS+RpXkU/lmsbRmSPx6f9/xqzarF8+0KgddQmJLlCLNa1GNDEo1CX
X8Jg2TIm6+eD2MComvLumYUspP5uu4J2u6WenAcirZAooB/AXEx0MhbKjJv66aK/
zDfbFIOu/OzSwOnM3yUecUTnR83lIO2bjZC4JGNo2uEz8A29PUAbWI6muOe9M01l
`protect END_PROTECTED
