`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ7VVl/X1iaOCQyb6w80J0vczjVZzR1jBZ1D3ZpJ/DWn
fsrHuk7pNecHFBVlWB7ELD/C//P1Bnlbn3vfdNHCPurtHpWgMFmucyO83AlrgZIl
YIGG9J2C+yNtaL7dEPP4sOI9BEu+UJD26vJDKFaTnmMrEVUrujiivHUACILnra/p
ZdkdupK8OeY4iGqQkpfajK+MXTuxH9HhnOtj1JciJX63Y0uVgd9O5oR3AGK2kU/s
+5O8Y5oxZ/+7kiCqvU++JkzR1BdhQQn0ic9JYN4pynPGC0mg9EDbisYnzyFl+HUn
njoqtYe/SaZeDtyTPN+2yM0gDgJvjLa9emP2/rvdApM5jR+gcd7N+8xWu+J8gLmi
eMpfHWrHGbc7FtgXR7lpOl1V++6TQxYdh9okOR9lHvScuiCDgYcelnbe1/4z3pSL
9acJ4Krn2MTZkk5Ke64vat74ct1NRYN2ULU519OuprDanBHvsVyjcISoEqiKRDQh
NA62o74J29lZZ7cWZf5OStwHIrXHrGPmsyWbgZt2LezGvxcYbXurrdgLXyqv1dGs
4QEF6N3ueH97kfgh6tnTtw==
`protect END_PROTECTED
