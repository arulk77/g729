`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/NGpj91Zthe00qSPWJbClSA/49TX1XlSTd8gvCiaPFxDyn45L8yq7Dz8oNXfkbUi
EvaHFJHhYuaOnzlGdlQk69lTiHEvYXcjIAWwOVHVAueA1BuPmf91Fg/16DgwMd6k
Fhn9S/P0V3kmYI8QJoGzL5ZDNfG+fk0jojnifhcybnfI46mqafqyVHapnc5245Ek
2QDW4qiaEFHDLt2xiH1+aWkVB7Lqdmyuqqf/MnXUQgLVX7qwaH+QwjN7le8vO0UA
9vmX8+hPJRRUKtMTK/fCj6kOTCkb/+GVzfBhN7w6zVdx3XLFns4aJ3Vu1L8gy82S
9UPDlNz3Fk2NKKadUn6UDRswtCX1Z64HC2Ivx8Lk2qBWDnvInm2JLzyAiet2I1YM
XhUt5YBSOfuJC4z0jdDQO4T5+yQxXrB79jaQBslO4H9srXBBaXDV87TmnbPlqPeP
Boq3o2NzHnZoW/9OAdKmKos6mb33IMWfF0r5L5wMDPIoPnS03H6uzIpmbTqrp11A
rKA3iueAc9XngD2v1tp7hTodYQ8z8C+8UWKoZ58PPXcvaodKHNxTSMnJsaCxDMQd
K617EZ+Xn1+2qHpJp4qcX4uygIj3vIin+ntiyc3dvfNIWegJOkv0D/lQ7fcE5ad4
OPOunnGcOq54eYYFUfogaeH8/F289xEYB85bFjS9hdE5eNpGqnXXhdBAwuE/oCQR
xIz1u9Q3pBgdMF3rWvSOWj8JfhuxwyXHC043KsTNvVe/BGwHglS7eumT98MVtTq3
DwxXwhrgBhfd0lacEfgUQRcj76Sixaav3JY2qabkDFjQnBiEqoupPG7GJZ2Y14NC
0T4pfwkLPurZog3BOymkJqUKlkWZv6oJMuCG8TgMbfT+6e5BCXoqRUwk2/c5TZoi
mq8n286/gmWN21zqJmyzbqHnw28J16a6icdur0ebGjlEFDPeJ2zN1b5jatEtmnBF
`protect END_PROTECTED
