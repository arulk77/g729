`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pqKpQvRbjNS1cfsuagGQ/BdxYEIvD8AQby57hvsN4BOu3o0TJpC54WSxCsZuHEqZ
yXMRSQ0ljTeiVrhOlWlz/tBVfeaq4e1kYavyLF4+MUuykFQIVxckvUHkgQnYeN90
shhxfnhLC2FQa9E7+sF8o3ekhbF+5EuMtCvPHrXTr0GqeZCZIfbpGLTTrPqz8q12
`protect END_PROTECTED
