`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu487HAypnLuOZ+t+6N8+5aadCceMQm5/fxIVbSwEXaN9a
Q1JmCKyI2VnT7N2vgUZC9WRoxFpSDYU68JJiB8gmSXYylvRXJdPlc0niqB1CFxuM
z9skeAgsp/6Fetr3vzYYWfnB+5McJSy9pYK44+Q8l7OoXtbMZU2HTgCHh/UFnZdW
4AE3SiHoJARqCIp3KOhIRzEFJssqMQKtadksyjObrc1sBPO+0TM4R02m+tOUbJJ1
2EMPaLqOeBNSI1WSfJnLZWRAf+gSFMascgvbgVMNUHgQpJX0RR2XA8UsGp3dk23g
qlour7ZWgkK3gImYv6oytVM50txrAQGBQQtUX2TvExTRyMtXKujd/gTLPTGyiIdS
8G1SU+TGl5s2yDIcaLEn2BxhcfztBC0f508554ljFRb8N4O9gXc7FdBW6sJ3FDAN
pAAgw71byFhH76K76dLjmg==
`protect END_PROTECTED
