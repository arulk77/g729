`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAF9xG3AllY7JjI9pLsFWLJDv8euPWqrTCmHFNaq300a
R+8WMs3SME7rgsv8g/ltpxqM5B71WDkUKBGvlt2Gl5y4dAglW2ur10uBev6oanMQ
JMtsLCVi+uRGiCRdoL/rhRs706RwHdd8fR8mDr+ojhxJIEYRNEzN2JnZoZPz+/C7
MVkspcHkDzYmJrC835UqWztKaerVcRBTpJ6VH94yFUWxrPQbGjRE3VoHBUhR4688
XXzWt4dXZcDaap7kPEHCxRCkjI2QjnbfIDV9MqE07YSBxTTe7/b+3d2bvFp7lv1C
7AQKoaj1fj+WRonogLj5katWJ3IktsGmKGLn1ESulImtgv3FUHg0cLOyXsQ0b9YG
b+yPJQdZvpdUBYm+iXRlK4uBZAKT9H5hI/9PEh4vWcZJa9ZdrfIRLXrtUp5KNsAq
sDGlPAWfAsRvsyw+A75qeRaFic4gClp7LUinANVyk7P+qn379U19xAfhPOQqbeH9
HwHYQkk8ofX3vCBoeielekX/0RPPVgfAgP6K9MyO5xsvqRXONJK27KdRXRw4V2+w
VMbK2D2YpPxX6GJ6YgBXZFM0HSaEqCOZdRYR5LJJ1XhjuFZkoiYH7+IW7PH+xlkN
4o+4ZKuOnZ3dowOdy0PqVE5mus7FQqE/e7/+qRnInfeL33ieCFDbTjvZk65M3S/F
oEiLzBkrjV+X36U28o2e1LeQNFUlcg3068RdK6+Ko5cn+7IQ9klGl1CrBZ7lJ5HO
UCOd7hH80WfUnpuLc9wXyEsRmgmWq82JS1NLt3wibNeihGWI/5meU5GV5Tvy4SFe
jDe7lVlbmB3PfeEVoDWoi2XgNUkC+eISip4tc/fucNYrl/OXsMyWjv5WKup/oPUM
Y2x8ji1GUQhhFv6sS6zVTtZ0Sic3XLJI+1LF7wSZsmCgA/nb34oGZDa44jLuRLMO
epgsEAZcVbRZI8TJOwh8I9orBhqMS7m36qbW7W+KRWHV6PS1hqqNqeABugJnn7J4
i2HDFDA5YrfOsyAXEZ/64bYQjhJht0RKilSL1q3PN/3/x9TqpzYgtKp7X8EGFvrU
ns4zN7eT0mmNrKEIGoOrvm14RVbJ/5+lq0p4yoFuVyMP8iunDYIXED1avePVziG9
aryLU8448lWK+KHF3majS3Y9ZsEU/pfxxdK8QHM9tu+Z8slFDcDauo5zvPsB7njO
ijxauiHrK97xMt5Cxa3JYdXtCPf6gRrOVjsmgAMkIhMLXcjAoISSqjHF+4ao3K5p
1Mj4gbnXTHFSbPSkb5KcCjnmEtZwPQ13MStF4sG/LrVB9cxuyuVV3eReibUsQ0Br
aa7br/ZjHwRtINHYJWQ+wUBtEk7nvjZhJEeomswB7fJ+hGVKzPxgGVjQM1sqe5q0
XhuGROcJTlVLnhv7vqE7/IqFa/9Dk9/+wKRgqyNcVjWpRU5kUC+DbcvoBeGclC1c
C/PX8Yoki1uE6HFch/nOgjy6ehfHcJYSV0np4zftIc8Cp06GbT7cYMw9H9m+23Fg
a0bI2IacDlsPcJjBe4KhrXYNG+f1IWkJuWzfH5SWbfOq637d0kq93EyvtpNmi6lj
o8/KsultzXpGXKV4ovF7/NBRkEEgZyQSg3iF89sxp7mNSR0zbhVl0rqimCywV6+k
BYuMxqH7Oyq15cx12J4CptBeJEzE8W8wtkOCQK6lxHkol8z74Y/w3pLfRQCExi+h
Niwd4D1LlEYpA61wbMYkIggX0rqI8QlUKFrfcJP5kR9LrLdWb/AqKW3SQJbmkHrU
0Ky7+4bi4QtTCdQda4UX6TAxTmMXeL6kJzhoRJar5XMKK7sa8K4QH5zspQ8/jwn7
JcbsKCAiNMgY4cXVo5ZU3xf7UtQXmku1CSn5AFs2n9i54trNozyd5dD2WGeWFn3w
Udcbh/TbX6i5QZmp72WEIBKfKs9LAMS1m2KVTvXN0iAKNV5m5vWcmcE6yJv5cpv+
om45NYA7HRycS6P9k7AlKGMnSMXw+OLyOPIFfF/bVDgBYTzsZ9lPPL60N8XU9se/
JIH6h2LN+SLQ075mThIXjdMuV1CVAHyuu5y01WHFQO/MZxAQCUpYzdDagCmwMzFN
215VxPvoSF/DDBPfxmzrsx9barF+NfYNTG9X9Jp/8mYriY6C8gWOusFU6FaEd6aS
csZ4nSKtTLgXbGQnQsB6+CgJ7kNA98YehkOLIQ9Qx9qCD5iCpeMdzdcIMys+io/O
bYVCoDXQ5Lxy5SIX94KwBoOummyIgwOlHduac/JUDXHZ/FvtYbzcWBPr98L0o9de
lQ/FAnpoNeXftAz0POq0ST2BAKqcXD57+r88CU2NB4b9siK9ZkoVF8cKidnXJsgR
HjFAj58LcXipivqlXZdIsYmZQ01scXULI7zi/cezbwHuLFvCM5V5s5S0ljygGCoI
mGAIwQFXsQYEwwvCCOYW2gMHlEHIyxcngndwnVaTFXBkXTLuJyMds7xH6xodn7cj
Eqdse6VTQVmHVL+JiOy3cft7tAbdmMQOQMNYFQ7H1LCsNNiFxHRx9VVbMpppre3i
BOAINIAzT81BShz2Dx706WnoiaIUbLCuWT7WVg1d4Ku+OC1oQ2uNdHB4dVgn1Zc0
MbN7usu7khAbGARnVnaPKt/Z0BEbioYkWuLrKlkuV2J14Y/3XOeNHG3vTyzxk59H
eYxc1QVxOnNObOu7XIkgf+nr0WRDLmV3kF5N0fYswroUJMvprwDIXnTnROTS6dj8
6ZbSLIwWkOD3GcOhXjFnyHEVsm7hGu1Q3QiQ9FRj6GXDGaXycWWRuLwP6fyEh5Oe
0lR6R86q7msfKkFttsSERNatndT7OeGsKRFzOiekWQpfY028vHTa0CO6hqNZ8pEu
xqoNeYALyCpPCZmNNKJdnC8Zxqf7Xu7RrasmkNIPN7lXGFI92w8OUylX5n7lDno2
Hu6Oc3/S7fcSC7G0M5Vohpi+mqv5w5VIDRC+HJXTmCNjUKaHupnatsBFTRVg5diu
UpodGWWH1eYGe73IpcJc3/8RE92/htEzZVVjvuOmthyxchuSbkCYiMoXki/3Zos4
nAc+Xby9hTHgcYWbN2mynMH1edY62aZmR4XZ+Zj5BfirzAd5Dq5O03EOkpR+JN9M
Lc5XmmZH6+yw8bMq4ljOU5XnC7+3/YsRTkZvqJ09bQ5S1P1RpYngFLcD/OvOoPyE
65Qk41+o/Pmm8Z11vZb1sSPEI4XEK6rRG17GdzlLAbZMKFVuzeoSPA0pUicgfTLA
1jpG5Kvgqhe4BxZl1MmI8JfXT33lcNf8+kBTRrF+i4DeElsxo9oEcnQToQb9PcMg
Y8oLxNdke6iMBcdZh69pCnSq2klBnz6p5lcXQw1JEpmIR1mkwYsQ51TBfOB+bEC+
yLOfZt0Nz0ApeH+ldan3ireLDhjZK5SKkB5hjm3AKzuw6YLq9FxpdM1+c2N4kLop
voeLBGrAdhzVppPVtRU2VIqR/jLKSj6xaxAG05NoZB9V9VtctVgSjzziYe3Twofb
CqIWBTHd4CSgaMOtyTLPFCBNCQA9VrbMO6LQfKowVCQ69s9O+ONz+Zsl7GflW7lm
eNDPej+n+QVikOgR+0uZ/PmK4G2XQasTxf0Kz9CCTeqOt5bfNFnLvsquZmJN003L
d5ikaxgL+J0o4LoXStH6ear5NJ0KD2l/zyde+vRrBUrNq4g0jCPVhyUnO1KRJFGB
nzkKz7UZrPlxR5j7JPHwECRqYjGYTm35o61YfxYAarB/7/u4I7kvD9qkSVpdqvF4
BeMbwruhrPBZSEZb+O5Aw0bQWRzmyfWu1qlBiO/dHTE6oRrwB6/6YndW2k3yZ+gO
W25Y03umyKhUfjQaQspRCyvxc0RrgtXUeLaJUL0ZEl8aR++eQrQosQQchda3Uxu+
ikSK/qM1yInMwGiIdqjpNaRHD7lR8OqDVwCH19yInUBsVQh68TXm5kSFpZHOGT7K
U3tR1mUs0rIrxIFGvdqOoswpb7fmm949SSZ9A8u9ylpJKYZOoA9qFJla6+WK5p3E
zWLfm+bdnjtAcjVMjTi2PGPiHtrAb5ri94dR9oz867Jn4Er8muAFtjHzvgUqaToL
09Xe6gVjZI6d8042jXTz5f8DPrT3ub2mKzhxihO36CNfBZbWty34mo9INDnCgoAX
jQnVIkRnCm1icV068nH4O++m3KzEo3Z/N29TBHFOCGrYRHO098abuUYuCosj9Cui
+plqJLNQLWvwj/qstKSk9oYPvCByeIDsUAod+h8gXq/v5saNxqd+Zx522zeurjam
OuLwMqLlzQbTPyENYB13DO844bADaPg31isMj5QhJ/cK4BEyKeFDLalF3LmiwlB/
pI3bcLXtWaqM/gAj4mekrFjHDgn+6/BuEh/TpOmn3pB+693832bK8LiClkCdY7i6
OWPQDqnRwL5VA6kYbwS1Hha60UadNiG6rJkNY46BTO78IwAGt2AcvR5z6dWtjVJW
wTyqGqJPVRmGfEs0sBDE28M5t5wn+kxkJsjzZWNNz+xf8DvAvm4cwk8vs3j3wAE1
/MJlwJAmCRGyVN64Y54z5WRrZykYrJtZRdkr+oYGfd1JwZQgs6hH5Q7dp8O0Wnk0
Kmb7ffpWwcp5HFjaALhzQp7e312DGcR79XtAYdvZ8wjk1hQFveEH6+n2azZZQfAx
72rrzvCFTzU6SPc256Ql7YP8sV5Fjg+9+NyHs18DSFV5UnCAiL82SAX7FOXBoIZ7
Nzfb4MMqeXt8AdZ8Aqek3MHPdqynNg8XNUCfDlIr0cD6pTWu/NINGS+v4MLxw9Qo
dM8IEIJg0rz/qRt+Oe+ZmyJ+v9Oj9SdArqGt20qa+cJvbbXODfT5Lp7vSd9urNhN
JvnR11iML06dFAmfr1sqUQwyCCrOfydXSiTq5VEWW/5XeDfPgqPdtYgvsa1OhMJR
nddxHgQgLNJ2SzzLkUgS73ntSWCsG2zJCj7SgfURCQmr7z3zct+oyiE77qzF7D2J
NYjJ9o4OthU1Alw6u/kFdR37netDgosu2arLgEQYLWCf2zwqgCyRDP5pWfpodIe1
hxAV8TM1TJ76dfYLfbGD1GnGcr/3/GhPL07yioIroMAD2Oji0iKx96fqY0pmIdV+
Pqgi9n1VwdSyS/jeiUkZ5J/1pKhmxkiXs2bkMNT2IZnTzP1mrU2ccZGiNdGeIRyo
aUrVwYlysA+r8lEjst7ZO7h22BYA09E7qWR5O2HE2lBtenhFFjE7INwFrhOutM9c
Caby4/5eiU9WBzxeSN9uBtLPcQzRW7VdGmuxcmvkQ5Q/VhkujWzQ5POTFBvU9zX5
6OgwQmDnJYkEu6y8wZBNAPDCnyuS/JtZkj6w2e36M3VmBDzDCvo+mHteNBmH67Mp
LXgtP4Wic2n/wfMV8aei/UjEsrj31o0gd9v2+eA4uUhKI9miygB2zxaBhhPuSIgX
i0IhpahomKXVLYJGMsZ9Aa1etZ1Qwj6CEfdBHxqe28/NyPvo+DlZMBqK9Q2UjTpn
kzT4FZ9KGVF5OkIZ13NEqQhlyQYwTQO7nFfi6on1erPGHTE+bS93O7RV9gH/Ss6X
TDj/du7xG7vkWGRCtGBjtYZmasvbHbrpHEemkY5EJAZbO1WQa+rZ9/RXzGinuV1T
ItOJX5x4mag0wmHw1304X8T8yspHHIWz/pX00vdrvSKhe3leRGwK05TtO9YuAs0B
uVNv9/HZI1gc3wy3+YqAB+DQyk17YKmv4QIKJEA3QbOCMIAE8cOrBupqdVFALYuU
wjoaXAu/kxX6r4zstpT4ulK+QAUiSwaRqKX5LhzXrQ0QfS1S8i+zySZwCfc4M/F4
iuRHpvuipVatekt17ENuGXHIT4QeynXtdaUBeu5lwRvFhu7wcrZTmEgwimv2Ibx+
UeUGEuT4Lfy4h7Et6enUEI3kJh6rGgObX+j5IaZ+X36C2KqnCjxsqk+th+RhgvGB
FJrzAD5wStblIW2gWRZS9IVnZrC5CeOlP1WOpGrlf3ygLdcGNYpr9pUVuFDH1bPZ
ivViuD6TsxVimVlFWLG0lPpdTxidwkKGCevJWqQ2Cn5wLYVSRNlQV5ra+itctagT
e2OO7GdZpEBVCDxsFb3bnn9KVDe6wTfu8uA0WdiRbxJ9LHFrdlrxFCdhiqSeXyXU
HqAkfTPNyJsO1GdQG72A0PCFy939krBrDiJIk/2PrTjUeQ5iv5S+CLmhcYLy8gGg
t2689LRMUG5V35BXTBSkFv2N+np76K/ye0G9aN/cccoJXPp0CcQZN8PD6L1Mjv4V
EyeDZyfM2MYrisPCF8eEJeUd1dCL8lGioOMOqQa1H31qR74DF2NjkkND7B5QbMSc
DjE1mHxzIr7IiHV7w6xo9Y37UPP/ckm2134836+dz440KcON67j7r3aRPR9d+mOM
nqhsIIJP1o3lNQO0yMQi3egZwttdI7rdVSQhgISt+tJ386jUSGcAIps1WpoYqVUN
ZNloZzXR0DWgjlqZFBhR+q1esvXSGGA6/quSF75SJf26eI/jrnNvUYSd9C5CohYq
1sc8DJk6QurDNO7dcSA8Hp9nJ6aImrTcDcRlJnDBHPqddS5AvLmOncCDTSa4DPyW
CDQ2gpXC6/QNz85Vea1WU5bvggZeC5VHfI+gyMyS/424KUZx+jcqLRjaCJGA0ViR
hrzMQHhEKDOR05PdaS21M/OSLjTOo2r4wVlM1LaeVLeZ8hQQaOjo9rVg0pZw+Jio
Ejizf3INa3LDBoi405etCfXfeFZ6cbGgy1cewfwMHFxrDsjHAwgUmUdAaJE/3AJ4
FjQXTIAuDNhyEDt3B2tYmfhpLOU9qdwpboup10l/EyrjnksgtBeOZlI7tws8LeFH
eHXr4ffrUQfUYa60CgVcN806IfDZgbhV3Ytwq6Zk/TbdFaibjTtWkM3zqJi9rZtL
fUQjWsm9AzKN3FHZROThBgv/4C6FFIsSTDg39gcBXhgl3vnlQqIlSE6HYXZQMyty
yEryizR7+narA7O6TrF8NtZpK1RHJeL2An/F8uVqwY6R5FBfDBK6i3xvuVUpVhQ1
sU45635X5nWjnPC7xlHeltW9il6OJLQ7WgR3ErR0KE3KeCa06lsszOwD1ayaJlwl
hD75RDeQ/Ux+eKFUONyiEBaD6Z4ZgGwxJEa+HlNW+Ek+vdHzn8OY/WDj1IV7ahRr
SCsAuR+Q1m5nZGA6xzJfTg/YM+58Jzk4P0jmr5RG923fVa27z5x5aAJdkfJSDVyw
eKoZW5NDspG6d2bJRIJX/I8JRBN1dRpQATVrmEkG5QIlshm8xCWVa/i5ieABWdia
Y6uAroKlJLzWFdLw0QZzaeRQ/jXUnqqWNKTP6//8X4TdskQPpLOLpAk1Qw/Sp09K
F5zX7whLiniabKrJTrxr8T2B/G5co1ay9zSuQAXAGF5IyE0hajGj4tEL8C0AeUbx
w1YEl0KU5Nca7c7LzMyVPLsdCN3LS9CGY0vSgdTIIyjKY6l5oR5YhiRmKOZhjucR
nahP/rtA6jg/zXah+QYMfQnX26rru9Dq+L2tPpu26GdsgTPZh+oHJQnVxfY1K1nl
4tRqV7n2bJSj554qe0S/DMIBThLF5gWq+fZeVvIMIaEwzMqm4FkoHm7b4VnQIU0B
nz3Kz0bKNtMxNWmtM9HiTLCD6ql2zTLmYA+/Nmz2Sd3MMPATqHVvxITvemHgDcRJ
BAd7z2t3mifHZCK4Fjn2B+bs4bpTJvmYkBa78DY4PRDX1HBsh8rjikYa/50JeFEz
VUJGR1AkNMcZjEtqN/0Bjs18eIxlbseCD8NRR0/sbaj56eokEMuT4GPZ2o9uoewo
m2LbOj4MTTKCAoYpmL/p2Lax4dLUNgxyutIBemuDhe46G6ltmsXJ72J6dLhuTQqt
7aJrUZF1uWftlBI2l5A3nttE0POu79Q7M58zOvXWJH0xeacN5bo2iCNAC4TROpn/
HOpAmPH18gebT6KVocx4Sj3K9Ts5tW9M/oYNAOPto8ANsY0w6MEjz4epB8bfhZqX
3vM+rhGGyvXMjP9camvmJMGNhdqf3kjqxXuAGTxm4wp2yoDY3/bqABJLhqJEkCWS
01y5ifM2g+khMP2/zAeW7LrWtaRBVFf+0Z+V9Uy5dhSgePPsF/9UJ1ufXMOdyfiv
9+MphTeWpgK6OoWdDMMWIHJCPXTzZToLEQoXlPNGIZStxkVnXPnwOAveZmypTJtF
nut3AVyhqKZxgFZaKH0BE8O1nB2oTPkGHgMkJz/o7gDtQswpzhz2uvAYt+S79SPp
Wz0Tf8xQlKmdbya3fm8QNfxMr6vxj5oeNGXhE4Gxe8OUUNiTtFvCqAvHtNt6J7Sl
1kH9z8NgclECEclQm2lENobGPSwXjUl4BKOPczpsYIdt7WB1/tkEvUnyJri9W9QJ
Xr/gCjSqGJCCFZQeAZAca1BABOmRcr7e5qKUlwsI5o9DtLG1bi18FPpGsZEshYdm
OewZgggbnVERcXf97VaVQL0xlNdKEV4rmTuMwqfGGUrExwe8vFbOEQvQgL4HwPe3
x5ibhRzVweJgmVqLr1hbxv+hj0x4C3jxPr49lXUGPqQ7XCDhqD3Md1MFSOvNYLAz
`protect END_PROTECTED
