`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKz/MrbIsJ66JyTCEVUxb7SqCAHJ+tfBIwQ3P9PeyZgG
wP9KPFWgecxSJWSWcevKgIR/TyPR0DZeWJ7t0SIPhUMKpOlqS1/Y1m/s/Zc0xiH+
JT5Tmy3/LPlIVc3OUgOQRxj8Ff75XNS82A1oEmzBhJG+Z4djg15L8xNFqPEcC0Fv
W9aLzOaGDiad8ANfj56q6VNSICqYK8pT2vqMZyl1L3D/lqePxW3PBSYD7x0BZurg
`protect END_PROTECTED
