`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePh6GIdYrkmXqNM4u6OvYixhFkU1PB5Erl99vr74wOXS
ZbeVUF3LYAS4L5q68pQndAnw9UcDrSD9rtsGzxbj+tD8cESRoXqFnWUbP0/M0ob9
uA/sXIrxLTd1vhRapZNJBZJkNb5yAy3LqXyqE8cDW5+8u7TkHuMRIsS3f+Wy5FnP
4R7t44EgXOJhVFgsvjF4zl5gwWW476UbB/XQr/nf0/ODB9kH6PLiQSfdkUj/V4+n
eo8LNy7j75C0eu2AuEHz3A0pTgRuiA5r1Bmwediij53UKCxJMn2OHigWC6XlzTNE
teVsbHFdFe8JiRMT72FryL6TOJOfl3tUqAfaoCS91qeMPx05qSHnFaOtrSAu0WJ0
BgOdjxkZEgNMIC31+H5KlHlMKMJJ6ITcOzVmNpI46wJ2bQE3/DTXXrsRecHRzyvf
iM7tYrsUYB0FhiPZ5cWxVg==
`protect END_PROTECTED
