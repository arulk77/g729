`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FztV3vTiecHZNSSFejEQBMU202Yl6KLNRX43qP/OKIlqUO6WEEsR9xYejjioTv/e
4/Ir6GLMXO8ZtuY7teNf33fHbNf6+tSFiKnvQjk75CsOkM6xgVdndmSkufqgHE2q
/LrObr7qLJReNHVjVeJkM9O5A/QElcaeFUtDIULsqhZeRWKsn5U+0QFWb5/qQ3pT
e+zPr9iIwd5WAf5j5NGoW1WSFEx8WsNKxxvz5krIwcyoktu1y0fLUgmcrZUhyZnC
GvlJ3ICdRrAAwh1FVxNsX1Zs/4DHFEM3VFFedRqI11H8En9lbPMiCo/D7T+Wk4iL
xyzhrKP2d6iyXw9RNOid3K//LXAJTMJZ+N4P4HwIjASp5Xyh8MTj2RNuu84hBf0H
bviAwmreDUmiKS8riHFGN0lMP674m3zKFHpZ/fnnCOJ8IMN+FkZkckzP6jHXLHYo
KixY/FSNvnXWxxDsO/O+z4XH77L2sQMih3zyi+fGvS0mci+D9DwTmfaw/mi5ZKgF
JsffHArEm2LuT99FBabKWq9LnYf1g+Tn5sGSJQlaH9AnEJsWTgbSoUx/MvVKoFzq
jkqe04+CeCB0bui1GQOmnesfttSTaSat4iO6kp/dA83oA3pv4TxLKSYp06rpSf6T
VbpwYDD4iISJui4u9eGObONh0h406rtRhJt+gyUbM/Cc9danUTcN8E/0btcyWTsp
6rWlCWIJQTv5PegHIiUhTG5z/fFul/tC36gYF5whIaUqIABkDtotAG1R7n3RDp/b
9Sgo3cicx1D5Wpxm7ZZdptXpXrWPSyJdrMC6TnrcBereRrwQ/P9knVLN/u1BmWN2
ewRKEMGSp4VeYQRWvffoUh7UYWUCC4n9hDOB5qG51FaFyYsLVQqQzsE/6mX42WL6
Vc26HYaZwKmUs5NzRIcYAebmMJS8p0WcACTb6tQIKtD3dIavdCCneey+Q12YVnbj
giKf0rHmIgmsAh59wnGtdlmQaEzp6BKxg6gh+rzlDitCUjOPFO4LQIAs6wdUTz/y
I1MF+2pNroY/uCJb1sd5AWn9h/D75dOdCiL80Z91ayqLttfyQT2QEEFqcwZPBNf0
3qOk8j8EGyzlUVNVhsW0FwM1myc5wtJqTlF43X1nWZU5uN6rKE1LqsdicGtcYBr0
ZnT7vYN4QGtXt7DkHu7n5F1YJHOw3ul8cPOOzpAPoD32ZDyVASPSv/a0Dh4BT/Fn
TTLX49twktcyLnDaFHAtlMqWBfCtYKwPxN9fptYmhQrDPTGwzroZbRhrFZCVXsu9
HOhWXPGY/tW8/tIMnznCSvsixVMDRUPz3plJ0iYBsGaY1uh4GW+B2JI/Doz8SJ2f
rXPeM24T2sddAaw46S9kAfD3MhMSJ57GdOf5Gvnho5LVAnK8wDuSsfUPlNDxHY5R
`protect END_PROTECTED
