`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZtJaV/VxPXNkSpY6rE5svPltd12/Uwy7cN73fMTPNSwVFFjhf7rg7tRtGLInx3ch
0o+18CEVWEHFXYRaviLfv3DwOXfb+ajFTY0SpfV+Y4HoH0Vbg9VzzT726SmbePTe
OByX0z8J9gSlLQqypulyIdIw+m9h44pCiw60cLfasDLIeCXihknpUyZb1wtudl5X
BvKCUz5aj0m3FffgmoK/5FFa4TzT4a1JuZCJBI6eV4HqJK50H5g6rSYlpMciNS7l
j09A+4xyg58lFJDk6xx77QE/Bczod7B0WsvYL3sHKzQ72RUdRx6mo4tVmjtSqOmt
YkXicBdsXPi/1wlyOkkTtN/x/ybzCNhD3KlXGtuiaek=
`protect END_PROTECTED
