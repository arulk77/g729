`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CxnvLjoSzUSiZK6doiDIs6au9c0Wow2u6mwvQ+v60FpH
t1hgcohWxBJyCWO5lGobGjZny1lnOX5v5uox5Tkt3Wr3MI3S7D3Yr8+lFTd8zJPw
Y9s8ZtcKWsomDojl2MXeXzaTv9C4N9pBOE6E4L1RXra6KexGg1edjZuhQF3P9JEY
rI4m/UjIDrOM1mlaqM4C5ghH+V+sCDZQ/eMkeWCOR0/d0HzrHfzPej5ADeVsea+2
CKWZ63iP0Msq8ip0T2x4uOjGwRxgO3sV2s8rfTfud/V5MzVDYLdn1auIZHWn7uGO
TvuW3rUEFbvpIJTMLeltgDhWzLHEYKryz2zpg/iyIQwhUdSCMidZ9b3gjiBWM1rz
BD/5RvBb1YpZE/1fYxgZVz83J4r+EivuLPE96/B0kCyTKsN46vLtAtJa4/dA5gmd
WSutyPoBYjlP+P6EepvJTMRcoyB1VlGkhLxXJACKNXkUZehwTTxw6ji48mdSGFd0
z2oxnOYVuqMfiVre8M9t0pFoJ8wkCL2dWLRb5Zo+O4mRXfex6WNk5LZ/Pt2Fg6GT
0pA0fJ4RazgClGz4gvCMAgpbfI0Tl6N6KWdzA28VEYk6bbb7ZXNQHGOB3mBO+h5X
KNJpO04/oO3rbLGHKQ2Dk9djuIxhmbXxOBizmtW2Mq+s4+A86MufJRAipdIY/deW
+Z1+wu8x7eU5Ia22QkL5aJhVcBI2ZHiAiGIN49PyUq47Nj8gUYYdnYKX15IIgDzz
GYKLz9NVRDgsoI3PWl98+UwRVEZZEkCARREg9Y3lXmKmXIWqeR7zDZWGYo2g1S/r
24El5RJ7v8dn0PLRkNTGBM2owN2aud+38KMQ6D54Z3hsfiTOeah7BzqOfjFkOyHz
xV0Wep6XbLWnIlo5JolecjS6QnSQfIgpzcSWE1du9gO6yEAKkTvLzoOaLuoI4vY6
kC3K9jV4a/2M7gzQJSpClh5L/uVpa/jadBetZFxXRsh0EswZ50Fm42Y3b+owCQkh
SQGtq3xwPz9BqaFePKqwUhnqQBGP8x+kfo9JXaOXOQmQmswVz7nCGUwtaV8EwUOq
FR+ZV8yKmvfweedWIBHwhMYaAQzYxbrXEutJDA631/KRYe3CoO05ym3GPE10a5S+
xffiZ3Y5r9vvsPLgW/KNH3Z2Uo/aSbzkqsQX45iwo0AGoB8kxISsli8yKCEXFqyc
jnKmJpTTqw6i+1e1UQuvnFwx62P47m+PVogaXnMIMYcwlLWTGWWbJA6PudVWRZI3
jJczttppkftB+vcr+jkEH6Q+lChQuxNyWf+2nVvHtRnHqJfnqMgPLsD50GBAgCRV
/E+YNl4W+USwnrFYC1NwIpwMjHhUnAd7N23dY/Ub1mvhZ6+VlHhbUGwE311X9fVD
+D1zSLyhPgdidAl5+LlBjrk7snjrt1hTc+76PuRKl8SN+naPyPYJrTPNZfFwkEa7
AmcoFrPzBhW9WxY3EiQZCQ/0EyVeh8fiQCkE+3ib7L5QleAhaDEmn+aAJzuFcTrY
BgnH0OZiLldDWd2Nm8qQXIQJYb3/bfFiFKaa13cg8EzV399cmQZSyJWpFCCutIj/
4ScsoKi+kFq5SSG9I/hs/C/HBIRgTuSJ3Bugd6yDqxKQ3HFzggefTNPqFGpdnd1r
GffZH655Jx5COOHuTCUyaDWmB7HPuoGeNvUtcMM3dPOtWx+o7eL+mWfYKZ5HAELC
A2cU3wceV5sb1uiyDk/t7U1YIIGmWMl9N+ckB8y6/E4+vMxQvkF6gZsj+muevzzv
Dp/UROPmOsS2ANoUwb3VMsqVoXY2/SpK+laxjuWzjTSSf+UEK7vja+eNyqMw5ImU
e7o/4ji74ZRGThV0eX13JO8D51k/C2gNSNUULM49MZtzHVAHLnK7jwO8wW0HDwdE
LKTcqk0v6h5gtCjbnX7Bkg3cD4KaGgVcKfo75KE5ModmbD3tgJ3IDVPFOfIPQVru
olWinfFyfYnAKAqPGjtNPTN/NiS80TTHKPFnMPu0sktyk4boAQ7mvWf2YdSfzTK1
mWQY55Z5R1LBSatxchYQqUJn6ZEjlQMnn2s0z+idI8DbQIqVTKZ+JBe4X3jyggCN
9YpnHlfHLj4cWQf8+tMuu4OATbRsRk79s/X2myxs9QV8dEnzvZcjvd5TrmkXlF3/
BD2k5lu2aEQySuoR9l4Tlc+x/Pffw22UVUfo26nz6wvCjWmnxnXkFxKIPgALJ9/3
oeY8xKm6E/FWIoryniNPsUPG64nQe+a6Bbo6r3z1soIyZSw5zxBUIzgLTuvAObYF
VtzRVaeMwafGpp0O/sY/xBOM1SF/LfHfenqTHHy83esSxpnRQt/HN9OlkQCHvTEr
3Tg0bJoC9yu/s4FxTI54ukjclFunHO4vTLdkE/cVLRoC90f3+1LFmMJpzDKIJDlP
HVbg+Sda90MwY8I8b+fq9cCwtbCmtEJ+HyqGmWuKbfLc5AQ0B6/c6+tbaomnx1hQ
s/hQxQVgSLEXwfejJJsPNMmFRJeUMeq3XqkYefbGB6EggDsG+t2m9FbptM8tfQlR
v6fQzJ9um7j2AF9mqSLpkYIP3QZYbsUYTneYzgqT5h1uio3am0cnAgE8+AoOb7hs
r0uq78oPsRrBrpN8lfIcxnvg3p8l11g3Ry911mTP1upLUegrebol2BuKmDqLh7Np
DuuyEfiUQZH9r/UXAWRaJV6TzKKY6wAP+/NHwW1H7/vNzhF60KRWOZ8gbBYQ9fy6
COkbbV6Hc+xNd2fs/Fy8DK41FDIYYap+xlJAdttRAoZQxTMYlTJPiZBBnDt64+bT
mnIh415IyJ//9evH/zIbJ0rJJwAd9NNAc7mW7nvlwiie1wIfF+3JltnEhpABNzF1
8+6LmiFdcbJ3liyNvcqoZWEF/17RQev17oKah0qUNMsio9PDvTvZZikVJFOUUN98
R/9uQdFPhxPcnp90BWYvCUAvgtULx/+aJhWn+Ueli0jXfHQi+Afwq6DA/rviBzXE
qmubBD5iaJCQU5YuN22HNGxYVa3tg1y/umqbX8yNjiixhqQAI/H36xvM2wJP7a5M
Up0ALHkULw0sxSm7KToMDC3N2aPeMWcp615n74jd/Te38mbefWZG4LjuIJLrA6xh
emUPbx4q4S+quSpnz+hcHAnCmTKqPCOdG+zDgSTt8kNA3qLHWqdagFFyweq1v6Xe
D2zu4N/k9oFNlnD79ELCNmvRN8L8upG0LOc7x/tdBT39hgb+bVbLV9Gh6UHqkKRg
UKfDi/KkdTY0kIZIHXjlEQ==
`protect END_PROTECTED
