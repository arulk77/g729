`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJODgcCTruncskI1ph4yaXU+DCxvdNrRrOzo3XApbl5U
XtInuZ7eSg0wBb8+K81Jrzav+oL7jHCiYlYgWeQ2E+440GZisQHodPYA/1yQczYo
OhFRO0DeVJvrnMwG3mOhXgBOpzuHprKrG8bTxKyZgfvWgDW42LlmHj60SzbMPEBH
dRPt24hjV2J3lgdhvSO+R8o3UhlD5DCsUzqnWQF6/UOHwJexZj8o1VzQJlbfWuAY
t+bFWA8p47OtxzGHX4Mt9MG168TQ+1pV+5+TeEjZ1AeJ8QWXh2QLkffmrNlurkYv
91JJ2RmgrRy2us2eTwA7DsFgNPu2zH3iL90RWiZe7SPb5VnIhNfzd0oPfJ8i0aHV
sFwbSLycbqJqCKk9zv0PkA==
`protect END_PROTECTED
