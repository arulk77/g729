`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yffaD8bntr/RxxRDyLVa2FtrdUzrXniVE93ZteVSgUI
2g/6ftxj7+lJX0sXFvIiIAMls9tT85qfzakGidVLpR1VPpMCQZhqkHRo9VNN4/ep
ZML5LjQDR5AHCciGeItpDWH8DY+nWgO8mOddsG8UUBKB7G62eKmZ44bnzlJnpAXZ
azKpcJoskmHUx1L6I2cpAiHG9HZXBUJ+8sQGxSZniOzP20KjBih1Jbau4KbVCV96
6U8nef+wsgOLLeHUFZ2prkmDfhgfxNulzw6hlk0uUfjhTHzAQo4d9siGsMalGuK6
HwIJRW7ZODYRKNPxLNHi92gkQSqHq2sPebMX7zOTd0S3OggKZxPY6pNAxhrZSOH/
MbdsXKN/1wKNcCzMtmve2JOEXoPbFd4PuFhAT81Rh8jiaspCJuIUDB0j1PDx7XYv
y4djRS3S2oGEJ3yTHO87wvlHcQ9RZY0d4ToDv9Pr0vqoePC6V3aoAlwiMnJlIAg9
`protect END_PROTECTED
