`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN9Wec4MEG1Xbg2dQ7LKxQVE0rBgbH/uoXaZlATPnrcm
TZdCwMHrl8EV5/oji0eRMvlRO03Epn3A2xQ8Ivd1reBRn5G0/17qoUGrE1991YjT
Eqb9HY7STm7YjxtFfjVERgbzSnuJCZUTj6QNO1QKClM1NlSnisGJAJj6Ub1TqEAC
tym5veNxDz4bmG/wFfM34sUS8YVtnly1VCkqwNSGQ+bsimOtOQrtyn9x/baDidtk
EnOwVtZfEgs0a6Sx99ikku1O8Qw4ne+wnKxRUIlcj3ez6YHWOQzrQu2IxHbQ6Zyp
2dIIYHUdWeKdfQB2iL1DuOZTRB/2wn2Xelc9fDve3gmBBWRvPGYuWD3FNUsRFCo5
`protect END_PROTECTED
