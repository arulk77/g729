`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
i18RHExlepW0j7tM2FzZzEzLz2HYd9/83MA3pM2he5sy5delPaXjyKTYeSZ6WyZV
aichq/IX+XshecY0Gzm4cnx0u8xxJEFLDK1EDNJuE/vl/KJP1C8xf3iHJyobxGE/
7+wicYsBsqvBX70Ol7ixrQkg7ObooAd0orHlMf0mmFpb0WQaB1D4sn9xqJuByO8j
tsmky1gNSzpo/BGpw+VEDpHFQ/G1Aj6kZ7Hgem7PTJYkxjf3KwRUGhK7NuBvIM0r
viHLL32yzFJnCZ+kvHYVCZSkYcBhQCka7RiVw83HqhR80YNe0l0BejFuqYvF7CIA
KU6RUyyHeTcGtu7oNw26eAnue4h9D8R4HT38G24gy0BfM7dhk+EYl4gxwbg4aK4M
DLZtGyAFTy5ABAQa9IYwVVECxeK20AFk2mGnvzVBPF9ERZyTOPSM/JJzJdihEjzA
P3Cfk7WGJWKxONttWoIKtKz0pGcHzUMHYu2f2MEVLTOEzsVH5Ky5wS8C5FkIlSA9
aqhaRWdjkoVmiXdXMqwRvOC4F8Ca2CEfLKNivSdLFIQc0eawMpwwPOJcg07duhmL
7MEV83j65BLdXqf8HiWB6H0adEesYAGv2K9Pgr0HT2THEzEUYLZQoEz2Gy+K1JUB
mb6nYpxPL1GM1oZ1G+6UNUyf3BiY/T1NdNM4ZFBxrEyulRQ/+TAupykTrgTMoM7a
uUafZWO0YE+AylqjxX3Im4D86ZTxiNxefQ9WLKa1kOM79Nlq1R7O/Oouwi9WT7UI
`protect END_PROTECTED
