`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIBsnDwYD8H0FWu5dA4GORZHzIuEgivIIoLOqIyHasdD
GatkPBqG5daO8z0hgmrmM5YqGpl6SkksB46e2f+HhKegh+Q5U9VHjywFtclpsv7+
LorNdktXEd/gMhLT0xL+aBihP1VMGFnUDtj1lulorcAoLT536lTx3shBLsIKyUpa
MdMMic5TmC7usDufNxVPLfZsPcr4RMRceK8HOcv00eeclW09iXPpDRM0PxrnCd9m
fjODm6vFoeb0M/zfeCrZfN7oiYiPeTWiV+VdVvdiZVVklyXAsHPNA4TLRPw4LSM9
V469iPtP8aLhwGLN9AZD+o14GihLD99osvTHZej+UrV2RzwGIBOjX9q3Crb13rOZ
`protect END_PROTECTED
