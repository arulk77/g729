`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SWdYt6eqZgdc1LqY8WupbMMGObvojOyGK288okNhUaL+
iKOdpGURMhcqOqUOdMryzMHtDa9ZQiSWpLb4gBL5PiqgJp6khey0zwZvNe+Vyj/H
KByOSZvvsFCm0/vOZleYsOLiEZ7GjxTfzE5qTfrbeaBJ9Abadba/fV9DFbevSTe6
ZULDgLPS3DBOkBUwp1iN8Yns70yZgpN95mvfE4C9AWQRKrbv553yvzvHfRN8iD6o
Oh+7efTX6XUxoXrK3LjD4oORr2qOmeHUVeNqDj/7lBKQIM72pLS2Bv8RSzZdphPK
kqG0XbI/1q50GG6V89J3z/Z0YazaQJy96eJzel44IkSsMO7W9XEIe+bREhbszT6x
JKoxzvXjZBVBUcm7ce6ZG3BZKcr/WgmAF982Yvf9r7Oo1YSvbFrMJ096Mw6vYxay
qMnz6US79NYGxH3JQax2bK5IgCc01+15mta0ORXkJHXbf5jhgM5G58G1KcdeeUQR
3fdQmcAbvpc4l0s8jqAJFG5rHlK5yMyfPkjefjYKmRSRuL68FAamIxhO7d2VL3DB
NAWTxwL+CHvzT/sIhLzloxfQqLI/VTTgTAU/KzGquLtISdbksq1WIrHwmQ8lKDa3
ce1j9BgG9gxwaV5njxCSV5W3al50ltwOauRIu5z0i+cHYu5xlvUGw9mmWImWyTRa
j8CeZB7COfGUxMn6Eg4Mfe1SZ9jZYdiqmeEItGD440WifglOrP3hHKTgMgz0MThq
jX/ttxrEIxcxzEOKWXb53J8EMqzEaMkka+qE/NJfLT1EBmh4jC16zQNfD1b+xtxS
BddmPfQXSrrSEtiVDM1DNcdiJ+ob0yDQV0iA6zTNxe3kqeHY8fsUbyVgcxVxcq5J
LP6HsQ9AexBeH5qTBR+0EHpDqokffILuwC59gu11A8XPNPBojuQmOquLiRs69rWE
JdfBZVv/nDA3wJZukKXL34sH+Degil4ku4QhPL3SVbL8taxHUwMZ04uTse7lIh4R
a9IVBJlu7j55aosZFEI8z5ClOVOYKXIEf0zLc/ICDeOq4AsdJqMCgFHxKMJAc19V
4bmEIvqAYDh6L6L+PXGLZyVlSOKzxC9X0BtYhOo0uVlo1XCNNiBuw3+72Kslgn+y
ToVnccL3A3Niti4oe4dQDvPdpuImu2JttcjTwDvefB7ydx6b3W/HfFBqUIoLwx9X
4dIAF26BUv9MtbynxRoFoxs7c/H+zYfY3KEYZoAhS5gbz+aLXcAIQoTpN9QXr0C/
3bxNvHiHqHH6Pc4PFSrmMhFNVQ0w2zvrvCvThPxGUtqo7OJ4GlFkgZPAm1fmJ7UD
y6FpuBkI5pIaBTdJGWfRTNbC1T2gt/ctAiAyU3HDBrHowRfFDC7o3ppOSA80U+nm
zB0RBiVKDqVYsDa5UAkZad/9/gBrcFYrDQF3W61GMxvM+qLhUE7jn5Iku0Trc0vl
UFLRt1z1+c6HO/YX9KFBGM27CaqWfiSMN8YW6XPCQL6Q3RITw3eP46Vu+8vI8tus
xAykAkgv8sVd2+OlAX4UNusTxFgwa/QKkWioSQP6RFMFGkNXkZ92jSqnYoZdgVuo
yoVyKCr+53zy/Hy0pt6TdB9QpnFRnEd7xaPqp23ibJa+fodLiaTkGzljGBRBBAD5
`protect END_PROTECTED
