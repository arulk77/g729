`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveColzmM835Oaknd2CmfPYF5fOvc/5UHhIAcPYT+jGv28
UqdE8uWzdGmhuMnYo8X6ITR0VTVsfjJfoA/114ZqlTCsHaD0Fy042csClMvg8/Jk
GyBQTkhVGZJgTUMMhMsIlncWl44d5DNSPk0x1OsMMmsGzxCDszc9CpR4y+GmYyXn
x1G0uXxcrHg/9SHyU+2MZ7dqMyp/HGyV7hPkpgiIYCJnXlB2CgfdUEzGobZsaWmD
YUflL0dkk8YXBKBf7grlaR2tm3iJCjEE/HIu393VKBqCZGicm7mq096Vs7Yd58kr
Dq+7qRCo4FLVDhJ3RPdbe+9eYSuRRmAmY97zV2DAE7iqBqj/B35cTgs0WJsAkRz2
9fHwo79aTd8cozhP4ZJQDg==
`protect END_PROTECTED
