`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHmTLGllgUXsnjc4HWE8FSkpVjnxtxtuXqkeBeIyQGqa
9LzzIe9rbQ0mi/ydobfjQfm58xd0NfijvA0AKJlU5OQmqSA/A+tmEV9Y5ogU1U8C
0sfugLiQ8VrYbcTj1mvJOgAzETg4mTeeIjG4tEcfChaJdxH2TCJRSJItZ+71P7Qk
8E4KBGRsntnrDXhnT6BlNUE7RDpEdNzjyT2PAT5WPrFgCQDyqIem6C2edJwWC1mp
`protect END_PROTECTED
