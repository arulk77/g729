`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePdBz4q2uzh61xVSU5l5Wj2Qmovdkdimsxp72ekZpgOm
PKSF6CulmoBlo/NbIG7BXzJik60Mx8rMpRORo3EtQ+UsvN9wSmRByDqVkiP9HEBR
YG2bumQs1lwpzitemHG9OZlKObk9nb3s/zpI2fA9BtjmlLFDmd3UI242UFlFuYPS
d6QjJRD8C4B2wM9gOJRApKVCkwYIfP1QUUW6roSk64D/cmOXbK6977G2nCTYr+Oc
6uAt4Km+6HTxaqEvhK3VFCJrCMaZCeWFFTP19XF4InVQDogdclifAM7iVk9LmO5Z
`protect END_PROTECTED
