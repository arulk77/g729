`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1acifvn+9uFDiG1E5aBW5XAi6JVbV7TGo8NF4lg+r/JCa
LN3ivPu+yfplIgYmUxI7YIIoLiyV1BaObA+UcCHFB9s7ib5uyUtuHR76LSYApgXb
JojRwzYo4CVnx9BIYsjoh65SDepoufYlz64yT5wUk/NFV5EDALdIPbvTljAbD+/e
rrWPNNvuqYnhW92K2SsmCWyxhEn3ivXv0v/o33SnOmBSQ3CHF7ZQeSbc53q3+Ydw
q8nnz/CMdB3pVvgZ89JSaUFqZZ0jkwOEbUhFnlsVohx7dkN27cgnQbAADMBZOpzF
JWBTPyLdXbsQcHiW8JlpTO93xvAcLKeNOGq/GaSeAwoJ5yl/3MVFg19oRei8hw29
D1yzFouwgC8U7gZAF2KB7R10ciubi+VGiCcidDxJAGSvoiuy61ayJISyqZwe8XG7
kI56er7BZsKYJWxMk4knVREBwbA+Cy4RkZd8F8/qFhsJXB4EOKeaJjTFlb8ZpiHf
fC83+SJ4cCbT8rSrQ91fX7M+YaGEbBYwugjVnI8RUTXackTvhzFDdkJVuDGcIhSy
/WBi+iWIBYoICYv3P7bioXuwh9Vnh6b1SnAiaHpE7tHTW8/gQMTbOZEmRzOOwum5
BE9mDP1VTy3BMMxpmqarfshU+Lg4Y1d0apiya4/PLMRbyHu03175u+0qhQ0GNzV/
`protect END_PROTECTED
