`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tFF0rH8vBm2htKu9WQhsSZrS8HQIpQmAAKhue47LSPpdbH+L/YTOplH8ApVycoNP
ae611nrIuh0wLqzFMwLdk+b9A2sE7DQTJbHOstq/AEtqB8nG8O9sHf/6TLjiuJyo
`protect END_PROTECTED
