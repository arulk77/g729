`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOSC3KPNQBo17HgVK0H/NU1R8pB+6jfxqVc1T51E4Q2D
CpmdAvma12/8Vre1nc/RKxxu8xfQluKPOjfPe9goCmw+YeBd4pjGfm0xQxBhCX58
KDaRZDtJtB2KUKTI39JE13IKfz+CrwhJ2+Bku1+ikWiDF0/KXfA4rhr46dyfoGj0
EnIFOPUW4GXeekO6qkCORV1/hMFbWyudMdaxgJ4HxNt0bw1Ls7Cjvno5Ff50vWdL
`protect END_PROTECTED
