`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePw11pC5h+mjGSFlM7T2fI/p6aQ58YKFaRGWsj/gkGAY
cTOUxCitBuPKqw24dnPVotz4yLR/DEyas60/fU9+BzR7q6UVZ5fOz/vBooAcxQHr
oV2igvPZC9JqzrfWe7ip1H39OzYwSZdB6OxPktlHFi0PjEoJzHAE43xhdHUFTeVy
/mfRbOt5aCAvO2HJxLRvwaGGLHvE9mM4UxQisPWVE+Zi1gGZ2hKblXOSyxd9wiyQ
6flNAS0k53R5kSlwRyg/hmmQZbe/Ysymk7EjRy5TYN+zJKbwGKnnICJtDe+8BT28
kMO4j2Hoa48PDjz0RMUI2w==
`protect END_PROTECTED
