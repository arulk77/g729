`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIObFoVIb+ip/6rfJ+f+k2A/z22bMT7cTzAmf1big7nm
74r/ZJhflfAnbnEzgT/U+PME2vda7LVETKJsF1Pgu/NdoyBadM3chIt+h82Jx8jA
ocgXXgbckOcJHa5CJtxW7ondxmTpbsfvNNIlJ72pIfjhIeog+1Fyu0iCEMHWVJ/z
HszkPybWfAvUGBkXpSE5pRd8S+8AwSUCgLIG3X4cXl++ov6SegtTFFKDGMTBsCGo
LB2QuC6UsMDH8m/7efQNWuc9fnCw8ciu7SBf2jOmquNCZ/ysQCQWb09P4b86TP6z
95tQIex/0oyCROTLfQhnVoN6o+9Eh8LctoUooRqJ1B+m44GMx+hszc8q/n/vsgJ8
SculXU54Wha1tE/J8M71eVMHqnyHecvlxV39sBA2gHFJqhssDOLjuooKbyVJBkpA
QR/V84zYBIAcJ9SLcaFZv9WSqyowTcyevXb/Q96M3nu5sB/hJzmefJAzUNjTfHCw
k8lYkAijvUedyJeA7s5cTu3JMKd2Wb1UCyrwkJFi0bmTfFmIebce920YkraMoToV
`protect END_PROTECTED
