`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNmShEB4mnA0hpuD1XieIzzwtWuE93clbJRsxcs7qouS
F1cPd6kHUvdtGbcyhY9ECl3hlIidvUXD4ylvW4AfKgBQtBDJQwOnxCDt/woX98sR
njcPIdumCgBFt7fIJMkTwI1dKC5PdbOUzDvwxH0SDzhLPJwJVO6lB9A7//Ij4iLh
0H8LFDLS5bvHn0DINXTBzsRMJ+3Uy75WhGMFJdQS7ZsA3wRmMfAoGJltucCqgCpw
JZlP76P1WLSMUnJn/ZShEy6RL32UUtAIvCuQ3lmK+OLIQb+482xi57a2FFZP68qq
ywgccf4mcMcuRXLpu+4oOg==
`protect END_PROTECTED
