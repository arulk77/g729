`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNOnBgqGdmmcsEl7VpBJBk8Ulc97WVnjLyGDQwbqeLVI
uFxUb0DepHFV7rBnqCu1QKColJvCCShl6Izk4/sZ0ZTP05OqmwCYD4mctu75lIUc
K/Q3eFABoQmgEoEI/lz7Z/FoWvbhXWnhEbb170LmrrxNIYXUk1S0Do3KT+VPzjVM
LslF3mHCT6hYaDOD8MGMYETAl1lXgrdCzoBULFKchlMok0vsvRuLh9irB8nnypny
TCnrbs5UeUeYDsX+BIjy+C9Z8SPZSBlm3tHqPg6uPdNIneiCZmptOSWcILLGElet
1h2cOAYXNU/0iw/C9hRALQ==
`protect END_PROTECTED
