`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN+FSfu7LeUsAuOXoJDUh2al2/3Xr5diILw67idRIK4fu
qna8qdjj9YoVaG60HPJGDrwxD9GjMtC+MDF2SDO4ryVQCc75m40D6vb3RSr10kGZ
BiSQo0YkLbpLhc1ALB8zruKao16HyLhjQeB7NNue0jelhULa4mca6r96t/f9tdrv
vRl0BPkWXz9BGEV3gYdezXz7xPouDqr3H10oV6DKifTgO9H8NSSuh1Vd/6Jt6mCd
XltBMX9MLMnUoyOGrO2B/09IGklIhwSw5IC1mx9J8AbAlw4usS11mon1BykxDGkc
n2kFIAANW6vBD5hnxDXyWWpoDjZIjLNcgeWSmmWJB6D9iSSSjomvNbM0iLZA8IKy
S0z0uWl+eEwed3z1Y/M7enDpy29UKbsNqFNdosf2u5RHpEvOHy2CR4l/QgGd8Opz
dGfgIWP0QuKQWnuzSG+mmiWaspMUrVJd3FKsIDtdUiPSImcbu9iv/1p3ZLNQFWbb
Kh1F/SH32dFR89cDnXHQp010sA4EakutLG4Ov67vNfmqgJs2xgP6VXYISsVGh12M
FLGiRqDprsZGgB87d9C23iaQgSC0oKCMlM5xsYx/vO4LqqLaanz2e2+XtUWkuonS
QoLdynaY99oknABi1ohyL05CR13rfoDk2OzYbdPR+/DVL6Uf5/QlOC9xR1t/SpWk
9ejdj+bgfT0cf27QGC/hPZ7RjxCYWU/ZqrhkFFyQ2rk5Kxa/EuBWCaJ3NZwCPu2X
Ff9gDkuO+oUeIkC4jZOccDmGIl5XYcgO+ZzxB/5g+z/6XSY+WH4dk3AfsvfY3oNl
VLaKK9dK8b3Smtw7KA8MYN6pEYV7HOXbLP1e78wsvfsmNhL/U80PNb9VL3uiXAUQ
Mco8FZxIqHt09mPeyuKXyVezwwtaPEZfzgzpaL1GZwY2f/Unst3odBeV6hL+p4v9
RVBqOW5avMyRDTaGfchH3BPkcfgbZ+Jimpxa5JuhwkJAmlUswqycFf5LJau/otu/
1KYZs+yJppghBc56hhffHNr5ULjRJhc6A8POL7NH30KPC+1+/lJfGhIP5Xl++wNk
gWB20l0wg6OqRf7J7pqJgabAV48ME47bCuA6GefVzMCdnflmi8BZWA67O5NoSxuE
0FmXuq8eCuESEoQ9i9R/TUNmeRjVCe6xB//uPIpErRnXxmNmhLFtOlTz74LPxlFH
DEiEfiDoyIhqO7JnRes45imMBGFbPoE1iWttBb0atZI+B9toTQYh5VOoRZ9IM/6D
Fo8WV6TN39gy+qbeXqMiUIpA8aOwdYSZg79CTPhGWg2xc5UQTrHm7EUc27sDoQXC
oJo0nhjcSFh4YJhFu0uDjTZ5gvPr13+KGw8Z8fk+QFIDmNN1+39EWhB+sXQIRDPt
wGNtUmWaVnKzbDGJZO2UE1vSd6Z613sYkNxMhhK+QQkcaSOfv46opvf2jZd8Tzz/
wCzhsmLxjAZxPVJc0kFcWTcRLPqxkXbueMS1xXvWqVfW+OJtyHREYz8uJ17HUW/l
MFTpfK01swdWz8W4fx1zEI9ugB+ZRNKjtrYSUndyDnmzsqK0ZYM3MGAQQZuZVgMH
DfJCIoiUsRZYoWHCrWk11PBYB3+imL6zRKlyWw40zaDvsSfl41CvUgmFgHKvdw3G
+4/Pi3WWu0sJL5rcB9qCfMzP0Rpj13s50FWFIjyTycpq5tJ6acS/8VrBMT+VBQ+6
IhCVIyKRnb9f28lpfNKHR671gmEfJ2wbQ3fh9YDPZOnw5GMgW/jWOyauOEgFYGhf
vxoP13l9KlhX8b7L5dlMgYv0RqdUUgzG2Pak3MR9ykpAcoxo+A++pZ3Mue60qQvf
i6xrIZT7VOMeA+Eykwhshx/FNkzDA6dLpPd28byH/yVMx67LDLW4Jl3CISNSO1TF
iNpc9or/VnVksDdrHfSzEkCbp4J2N897ncrxAcFfFnKE/d2ypy40B+bPg5dXEiIi
dxXdPJS2NjENKwMwu+GFuVBSVEB5oh2dH0krGF/uQo2NtS922e3W0hoQtD/9T9xv
z0kiXiALZcFnfhqtx4YgipeFq5AY/rynktDmeKdplLSelI7Nyhbq5cl/+PSgqQb0
QdCEnsr06t9IE0vkTBl/6Xvjts0YPlihl8GYn5ZO5NDToG5nx+9vOkuF5G8Yz4JQ
hhBi3cfW6Yr6mpHF5g0RZuW7k2agQ3ad9kY7ebNJ8HTrCxzwwAVsXE/uCBfgjQYI
UTvoOIclrmd9k79R8R1brmLUK/TNvL5+ZDBhdjygrifWOsEI4ojIxYSIM+Fkz57/
Rv+SPuv5rjuPbsrkfSAq626tKVXspBZCnFIyVggmvV7K2azTmO7gLOR06JEsfeMX
oYoVY8iAroSFTGn4SXu4HWwG5hHcZgtG30/9V61Z1VnGb6iVzJ6ZXfCqTNq0o/gA
hHE+mY91j3t/TT4iZPVYyk2i7U/Cv+YxGJKFZjTBPmyRgbquJF7neCKAeX20Cszs
/1WxVGh/qQW4Sh2xmWcZPxK0+CtA/T9YS60fZFZt73Nly2VxHsvoCSgNLu8v7j00
v/uGZZ/dXCUkfBRPYKjPtbVfO/OEmDzON8msIt0DeToKY6+lO8Lkdua9PayjzbWj
rs/GjqRqeAFLiqcXoa6GaAKmIVCiiXa2zVonjWgHF1rKjufc6/YqfYiQLobZMKYR
a6SsoXp5IKv/ztck6M3XziMDtPGQE8eRRZ4k/yuLIPUT5kAhTaquU+JP7qDzJ9nG
tBQBjjHzr4XhOzhaDwxrRLF2skEpWbgFRDz+7Nk1s3O1Ihdiglu1uHtMmXJbIXnj
zHuPC9YoT0fkbZFSosCWL7wGoY9mnX1+vjIbrvsV58+UWDeamO+ZBWrk5blwfvn1
OGxncXL8OFiQavAXopz9/e3+io6Zwn17pdp1wToOOUKbLuNia0Vf4JsOtIt+JYn+
LcyMnwngxJrgxAl+7nzB/aJ8mZUIwplz6XYDgvjEa6uynf7uZp1aP2fZDGScp21Q
/XrRUyVxqlcCwYzmBDAuB+5qF+zYf1XIMkxB3VjU2sw=
`protect END_PROTECTED
