`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
yYjQ7IPFihZCBc90L5yXnZMySLVrNw2Ao31G4MGtf14UIO4Z7Ki/tCs6GPLv7hdE
vynDgFJ9AIuwJP4eqJg7FYhOPvFMUaPq1Djsjv4b1xQtgKYhdZ8meVQbgNtvF/0c
P8SXQhqQ4C0RosvctpsKWokH/BnQxGKQIQ2jUHdjkxPmn4MxuWawwWk3YpwCZXcN
LnKnYGlW3dbHQ6437pTtalzWbbOh0AV3kbBVm4ulEr6ds0b2NbWrW+zawEGVgjpa
J+CIfSPzXFfHjzq1EswapcYG0aPldv9HbNtUHYWm39dycjqaXi+UC1REB/xQ4ISH
fuBFjiYdmctBSy6HPcSMzW2TvYY6tQzeC98wy3AcsXIgv9awSJWbXZ3fEQ9OXXqw
K3+TL4Xobqp7MdVRePX1DChKMXijKX15AVJYT/cbaSy7zwgcyKL6XZv+hcRyjvMy
MZFU4F3+tabM5FH4XAfjzDp8VD4giqYuOcziTp/Ay2EcdznUtFnthjdn1DjPPSJ7
ZieMxuttQw6yxKxjtOUfUBTstAAcZCQL7egLxsHgps446jQRqFiN0v+4Uqr0OW8a
4rtzBGf/TErJe1kgnbIqilfm6CpoviNyeNFFeYZGDNc7fiQdFNrIQkLcI2IpyNQ4
Gb/iq/nt94KD+JlT0puzM76cZtFcQQihksCPH1C3crWXLbhqdRA7BwNOSDgC1s0O
1mSvGpuhwW2KTi3ZY3cz1jhEcP4ZwV5f1AusgJSz1+KCS3T0SDmdsgY5ChtOgMk8
`protect END_PROTECTED
