`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHgAlQx9xOPp7U/Drg8HTGVNFHPTOiunN6bg50K0HX1X
2npcnE37Iloxjn+MVcTPBLdR4fuW6gQlHLfJuDkIr9hBZRl994FwIOyjIKZ5Apxh
dAuwtK1CxvVoPopTwXt19M/uZSs2MuLEl0AWJbN4BxLo9TDMwTDdYUCbZzZRs6IB
zWhwVe7w/oEY9To5poT2zJOPvvPfG7+cRCSj5CMbJnyaxtj/o078CJQKNc61kRKg
`protect END_PROTECTED
