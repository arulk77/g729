`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48G4Z9C4QAc5XEr9qFe8YkHKckZvqqsqCWEauvN0nB2X
BQptMkmKs2vwfFuUQ6fja+kbT+H4VgvWSFPQ3ZEPCR6Z7RxaMpEp4Iif98lHGWbp
LDLWutuKI739VO6sguLjVbcKrwoK/4c0LWSk7urDhciJdL9hPuQ91IAGuD0dp85o
mlQUeyRm3aOd4hCRdfivbXe0FVIuPOPxzZIFCcQko6FhM+FiCAEj9+gnZuEhCWHd
oqdL0AJ3axQ2YYY8kxseRMJGSZrbCtA7RQQPT+0AMik2qcqt+NpKKLSZJdKXH6Cx
f27N++++HEwulAt45UO8kgQDFFo0B3gQfR1jzksYFhdgMwMEn+9pLxG+lPW3vqa4
0llmoSu0CTaFl+JqvikWG+q2kfftFgVHJ/Nc7A57Jr0MrIcJpNAAt/QWF1Zg+K1E
Cv84tTdZoLLiFW448bJzKmCI033rPHvzxcPbbKnfGhVhqt6N280/OI3JEA8yR76i
`protect END_PROTECTED
