`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD+wCXknnL/kg2NVNb+94iCCPKl4mrAAd1RBD4EbEhQf
2oKZLC9PxbG/E0azl9iIjXtT7CfsOVNdjeW1+k5Qn+Bm89A2PA+YIkqZCQ/DhZJc
rNHb/pfwjWfPcQTBwn3+k2bgfA1P0vR8pz5kq0YXx1t74Pl2Bf+KQccguJ0i6FQy
kBwqRng2nqcdhZZ57CJqm1uHADSSf2g8x40q6DH4XycYEhr7bv6iI/EuGuiwWk9P
6eeXhmiSbCfC1SFZmvlq8pFe25NAZ4b56F0UsSyStVwwnY1yQl6zllDiH8jbtNoI
ZYeGYkbLQwDbRTQtFa51n3pT8oPQXifXsMl8PwNp/Eq8BZdjF0Bz/tN4JeZDmSkc
SQ5kZky5C21rAljD8qzvywkzwYA1o/3a+WYZ6C2w/216VoFPwY16+v2BfkSXB8Bs
JdvZtQHWX4kw+sYGhyuZDQ==
`protect END_PROTECTED
