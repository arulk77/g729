`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN4OVVinsBVOtttXiApitlVYm9ROkfCq1Dld5I/82nAOY
fDdCk0tAgf91bJJjAXLq4FgM4oaZKjbonjfxT49jhY9rsPLXvGU5b0RlTvUmd7iZ
6EYWLntUXTZKQHTMhMPLtSNwvWSSxHLWiBmrBkFUn8gkVL1bgryA5VIbs7K6vpzW
v/GUjLKSaTCEkHLCVBQohwILRnAqVg7bxCt5Vplhm3YG2GN9Zkjb6q7jsZSs58t+
5JkH7y0tEDT10RITIR6ggidW49DNCn1kzY0nQhSWKCgitJmJNDSbcPCz1CjW3Ezn
k2TRcuRP5qOZpN/zlyXSng==
`protect END_PROTECTED
