`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0BzKPAl3AykiS7Qs/eyyRnO8Y2awsFT9VX/OBu7H59496JTg3aCMdH8WXwfYjHqX
BMQqYYuMq2MYMXOwiPsllVkZCETwaKmMvyD51wAuNHUuFg+px41xSFwFLat5lI1w
nspBIZ7yTgzyMsQb+p8RXvvm/GgMyvx6uKgHLgwFO1O38+ukzo/rTwHW0ZXQ3ZPd
GomVR/SJ1jbZ84I/MABmMf1R7U1Z3hnoLffHslZwEAD9lIgGyF9t9OODk6B9lnuS
Qu2I7D+l9nSnHNHWdBCNYzHLQ2OaVpuu53QhhXFVZZypnw0FpXFJ4oeBlIa/jKIO
XGzuyP31sXNXSaOig6NthOhr5OWYKC+i/dXM/RNfXAR6xxVHRygOk8BqzkgQBfpd
7hKcQ7Jn93ytum6cDqh/FiQ7jXUQ7aU1WTJL+pzR7v6y6VYUPFKg90W9w7AcQo+t
7fJTJQCLNBb/lVN0If47SKD1pvD6Rybqrk9+iIkKRRWK88AuYs0hSCqRNVc8/OSX
JaRIsDn7Rfaql2n+bS5bMCNXyyOyFotVYUprTrqef6wbn806KrXaXgrI2xc3MxkZ
R+wukWPy7zH3gsugZQNLH3gpJEdDOj+sWunY/r8yF2oEmqe9VkZ55GyEvaro+s8a
OriItX1Y6VkKrg5bLtuaFiDLRPinXmCeQym0WkqFH2nOU13xrgmisMRK3238LFXs
6FUF5WUxKatYJ1NvpMqRfLidU+gmYHjhmCU90U4mMXktHXZq+wB5hlX4jbnbBS28
jaGk3YX06L+5J8NIf9YvNpM32vuOOGhVa9a5AZAqOFU9Xqz2xfTv2KLLKQeejSEl
F/pJd4rUORp9vRjCnajgzoL6Jl1O42hy+FjLlhUS+D05EKHFLNBiXKDMw6dRP/WW
RIo8Al5lC+Qh+ZgK26MvlCUbomu1Y6y6TRZ2+uyKNLuMHnpUteQU+0imakeEyjic
vT/50qci5parl/bwW3mnew/XqE0lCRv/xr1f3mo6BkhsjSPx0xxswqsTnaTOLkxi
IjnRPClr9MvyFys2aYG0V1m+oOgA2yQFioY6ADM6Qwlc2poiyCsvdsvc4bufurmo
Y5AoP+1xkvNJ5qzFQgGeO5HiD8ajFHoT4BfqmPr+8jRC6cTsKMaY5SS9XYA/jP9b
pt6ELTR/H9tZOb7Kn9pxP6uUtLzRMeZBAbp2wsI0NtGh8G4i8Ujx8w7MBw+eAhx2
VtXcLdKy8h6R2W/5CJhmFNWwEiWOcxg0SEIcTqa65Lbmnn7/wHLtWd/ZJc/CfBJp
3HFSNS/pAJZcM5ZiMJJ6biZHjSq39BdqtDgQsWprTmaS1mKBkEVoc9ufhz6s2PIe
/KUMoLYpz1Jtqd6l4BbeudCVKVHrdrPO3YkNE9s7tT3ThI9NmbY0/Z7OEOxUFnWF
PaqPbu8/NI6PLiJKn5lL9XHAtcDakRpvXzocB+LhDORSSdtZPL/oUTkqPJV3Qv7T
wlNYFv2KsqScnSTNbU/DVdPUZYgSYq+SunbArV/Y+dpMTW/1us/JTELl8FIMiG/D
SsdqCPI/3oekf75BhKKAoVexR+3O7+E3qWCZ5JojwDA0oG3qg0ADAzkh07euG4TH
T2kR97eVi4lBU0pE5ldMOOi4e6zaWKGttJMTY+qg9mfQw2X2tCSXYSWL2ZjZ34vA
`protect END_PROTECTED
