`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
EFnFEobTzADQey9vjo/iB1M9TgPQrbGAk+QlLxDG+0JxJPH8YT4uoKM3NriAtYuA
k6V2x0xxFwqjb6w/gxAbFczm8k7iVM0jVmDRKwnTK/I0E20w3QyyY6+6cs2CZTDM
KSBxiO4h5YOEsQLNH++TVP5Ea6813KN6S7em76SVY8xhjxn3XvYM3OtA4oWBLhK4
`protect END_PROTECTED
