`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCKHNjPLiapzF76OXhXQByNfBh8S2DoF9NcB7vjxcRUJ
QT9S2CojRaCyMF2A+Lg/7XxBD0LjDK8ZlcDexMyk1N6icqBpJUFkdvEDfQMGaQ01
nwItTwWY9Gxp1ausUUODBKpCv8sa8covIRiSaS5bj2C8HJvmKUMWc0xPACgvXzn0
6/q1fEvm0Gkhhm7sxHc4UXLIwy7g3Edjj2eGO3bInqhuSQZ9DQVqGlotyU89Kbb6
U7TagfE3/qbuuAjJBxCd880L+rjoJ9X6YPI57+b+t6jD69jhAPvs7fA1c510O+70
4lajoyVanmKnG1/0urnh9K+9JQkwJqQX1o7faNE8yL35OZXpz16ldLLs02HQXM4F
tND0aXn8pppGjitf0vbyFkUc1FrxIktSOG20GR5y0AuvtVNyWArBG9Suwd8uSbri
zi2LF+EgXYVbPnHWaOze6p5QOV7tThvQMRaGjpf2QKVJ4xxJ9jA4Y54hVbCkAjtV
JWT+Dzu6xMhAhQTNbBO2nkY9BVZwkE0UpaTrh1MdWlMGS3wTAwtUFYFd5Es1xEuh
`protect END_PROTECTED
