`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIbcFlUHP6n+AkqTtLjZRhvl4d69pEEE2iIRbIHNJ+f/
t6DGpHaHlNc0sTvxLGII3HP5dgEHMDMMFNDH9dgpr8MzSBvQHu1c4gRFXvck7nLC
1MbVVHsv/vNEGVrJYPaaCrell/HO2ZBaOpW2hdFU9/0ID2NrELLT1hVK5cbjbW5Y
wp3iFtWjw6nUTBWq4X7T9vpDMcGRrI5AhYRa3CD21BUnYLwbJ6qlnegFmWPH0Ssy
mhEWsgQWGqSlBplhLCSJ4YGJihKl6nash4LvceoES9p8A1ffOKkMU7CpEOLOg298
EwtBb/aaCvWtRlyXROBaPQ==
`protect END_PROTECTED
