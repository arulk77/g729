`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHoQe7h74VxmQ92ToY3ybxil0mRCAOHqzVfOdqCd2y2S
rjCQrRFU6qgHzbBVNi8Yokw3C+1kqFN5aL8xJNVBLHtr8IPnjCAutnUhz44oI6Ex
vka2csHNUKrqlkFCcacLUOMq2biY8CFwcceuuC3+NvHY59eJKtIJCGYT/nnjajPW
IdvqlSq1RaF24uRrXhJg+6MCh9k2/9LYIevCypNFopyowWxrWRBFjZU7flZdvYNC
`protect END_PROTECTED
