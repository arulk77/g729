`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDpxMZmwOyQecEUV3IICeqMa4Pr/BJZi1sYDxdhzltIm
tZDAutO37YBNGM4KtLk4S1Y/XcJo3NYbPGOM/gWELzwTt6UaLoBNxH2z+8V1G2c3
1wRl6erbYywbwboj9G1jTVsViwnk78UQPkIuZ+9AJ4k4J4090F4WLUAurwBVbyou
L1Dg2b7irQVVBtNO0ktqVg==
`protect END_PROTECTED
