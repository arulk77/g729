`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4x/d/J7fwxBdVxVs6DxKwaRQ60PblSDeIMaxXevcvWp+
CqMHED2g2XXP3HWaZxbNanCQFgQRHFttTqiAXlsg5EHq09Vg/qa6y0rse9sQO8Sz
dNOMmnbY3THyxBxHIiePnSd+6vZy0NEiB/R6sumvyzxfbphGGGtmSqxnhMIqAQZa
AlBqvII0cbqBxmQo27wHeHYABOLgORsH3LcXvnf5oO9SDShV/d/bbeypSX3WFRx/
jWkv/ypR5yzUj4XRYFJLOEcgCnnSPzkpV7PbewUrVw4=
`protect END_PROTECTED
