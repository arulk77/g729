`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIYwHsOYlecqSilIBHrC08znYJsBpeKq5UU8xA97QUOs
5S6bnlvpaW/YjpPflMqscnc68yt4CitvfXH9zAfbC3iPi4XZRQOjCYkjoP7QD004
eta9S/D7PHoD9HP6Ds0W3n6dTCNS9Jg2Ca2UHMjwHjMVsEa6pR3up7JbBSYTfYIj
Ef4fdcWLNXpLK6QawE8iPyL4mGunlLyajyaHNc/IobJgf4F4i7yPfbUuHcLN3XqY
uk/aylesKAzD+l6jhzglLLBUtjousGjAZauLdm3Q+oMq1WBr47F8rTNf8+sv5yrF
ZWVnjyRn2INSvOQTsPVb/UFZn8Fhxp2FJ0o5Q6dr/hfeLrDgOLFtPdNru4n7HmuV
CPA+JsX7RaLzaCI7EsllvA==
`protect END_PROTECTED
