`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF2a5l5LGmCL7ofJoU9jJwWJSu7Euo8A3WsflPoFsWMz
P3TOA7404U8hBI4DDQwsZ1bxt8ZeDN7w/0Zv5hM5IoXVPt8O6UFyhSKalUStCKL3
d7eTEpMeOu+/A732hcXErobaPHMwJg7sG7/mgXJF5bf8RL8LKLX2bXbhUdQX0SGx
wS43VyCf9wftrPObBOb4c6Q+c0ZR53gj5nlvql+FmShD249Y1nRMD3mup3xyYGUe
03iyDh/6Hqhpa7OeRAn55RPAefS23MTgTVv44aRqecF1TlkrGVboip1eQCiunt3X
piHccIfKi4qi4L7UqZlRMA==
`protect END_PROTECTED
