`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9CNbNg57i+nZzveqWSPFbAMeDP+n/Y9bkjh+Z6sOqSCV
21AOtb4GV/fNKMMPn59Yjcv6NqMjV7kjd+QtWc8B2qESNHQvwSET6Zz/Z0GENhdz
QlmlDZfPCoSFDaPftenEKuQBSV/zlJTx+DgfLFOc1wEJJ825ucoQ/himQD9kkAeu
lXrOm6IUZ18v8ulA0qS++oa8htLaYpbQzL+o+jPDXWX2D0g0MQ61ni4eTAhy60BL
vZN0OrAu7fPjRDvJbXcxHhP2Q4tDkJYAtEOQygMQp86K+AUN4WGzhipvjxSruuqJ
sHXomwYewuz9uX/1a0mnwaSEaI1UfE6RT8y5gmKM3Vh9yTRDEWvAB9V5l9wwhTtJ
j2YIZgcmpfRiVj0KAlC2GK4k7RIvowWX5KLJ/hQ8T/3vNJruq1edFx+O0HgEkDcM
Zrt3M9f8N4AwM4RrpOVw/b2g2w18ErV7CBY3nY0fFeA=
`protect END_PROTECTED
