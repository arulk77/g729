`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C2kEdzI6iPi01IPM1RAv5Q9NLLsKFlmtsK1yyqq26z7z
wtuYFExZihkxZ8cBZf8+cc1wIJMd1UoCx/JPr99BsjnYriJh7RzdzK91DzY7sYqG
1ErFokyJAYuDo7lmuxwl9YbrHYX58uhTtvU2cuMKDH6ZAkI21aQIHce9Qp021OPL
ZP3U6bQu1fLn8Z0Fk3gDSHujhWvHsurLsDQDnIITSkrS0QQeBgg7aGGu1jJkYz/y
f8wzT48PJczgTHzsggTXrfi8mPOXoAGZk/QIOIiWaclgFag16a0ZX/FaKMIA4jHX
vb4ougxUAOHRkZs2XIApVF4XooJW/Zx30s7tmL4hRDuB13FxyqLALpT7h35Ykp3P
WS426i/fBZEm6HEBtQgNVugMxyzbshBTQ4y5he+gFapfxmbqobnEPBUwt5CDhMUb
5KCcVkfLnnMeqYlg/HH+MEmAgf4GbFDIFXLaD4bkeF2+q/NfUfcUG9dZgZAWxpQ1
kEsYDkfCC6BLRTonCrT7uFrAIDYECoedzOlvRfgfB4DYti+o2+Dn1uDQb8yHwWfR
EUGoQUJyisDp0Ns+qpcxiGRiDRDQz1c9mNeNv8C7Z77QvVg9ezpAtUovZIbs82PF
K7vF9xQhfkm90tEkAIxFNhUBNLJ92OI+gvhU41hZzrzqeRJDrpUG04FVErHUdOFB
EgICq8VE3nke06apDkWTSDiQtz9Y6UOzPwPXpEW84qWS4j2iuYlh8Et9Dp42ejQk
b+X6KGpAoqGnJOfJhXh8T2Ij40PAHUfEYCdZdn/07+ZR7ynQFJnIwiQyNksWLh0d
retyPsNpKi4sZJwC9IoFfqG/OQ6gI1e/VYKvK3BjJ9R2y6gIfSGcJxlGhc5RrMKG
`protect END_PROTECTED
