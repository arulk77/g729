`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43gL1Qq46ZYZ5kcHKbKRjoP1nz+WvGqZTz/5zIS9YjZg
BrP6jom5AKe7RcyEc6RBNaFKF9R52S1B2FdsfYa3AvCdJg9PAxvTHfcG3BHci8hI
CgYoJsdTR1d46FouiYg9sbClvwfh5zUT8rSlnfQeAC0=
`protect END_PROTECTED
