`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
w+I26tDvvbnnvF5p1D4Ko8wil+27lnVgzbAW6DIMmg485CUcm4r1v19JrVbW7ahP
/qe2UvDl+nL2+WIUFLeD4/TebCbZe7Z3845DiFVBP06zJzseCxQ/UTv7aTaGRwz4
uzCERA385flgag0XTLMkNlDxS9h2g9Xw+Dqs4paYug79/Mah55A088W3Rr9aJd6r
0PphZ1zwc3tuJh2Ss92nLgNIZJ5KZ7AaSF+KATMbHOo7FL+mzWv0RzuxoTk996xd
bHZeXu7t/WxLmtWAcgSP6O1DPwVj7GpQI4mtTawBHk6llSHGdVTjyzpMnPWxOCza
Fy/1+s7iN0LIZwX/6iB/s/F3hwWSwfW9q8+CRvRr4Uo=
`protect END_PROTECTED
