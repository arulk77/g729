`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLF0gHiZidQG1ZujTmHMgKqsAUqo//E4sFDh9Hs5rppl
SZ74g6Qhgo9sZT4m0Ii00pEXAKQOflPJ1zMLk6KDZBImx8TW30EyL5rMn7rUI0wA
W6vcJqr6h2tYkrRA8iPrgZAD7jHvbUb2VZZyFalzjAwYGOqiDtdzfUdtb7aaXyOD
2FCMSgkzBWU0LOpsQOQXjOs5ntYliKU2TzPZgyPVGLTei/XsSJoMphpLYu8sP7DH
FHgoUQyQv9wgQtR0nb/DM5MfCx2YIzkRN5Tb95CTz/rVqU6MGP63cV6hJ3D84Y5t
0jhJ6fRFC7G2ptYj5v5pZg==
`protect END_PROTECTED
