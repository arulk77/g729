`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMFktH4ouUKV8y/HLvREh9vJyp5okpEItosZoMR1Q7XKs
xIj8sqqeOdO8/I8DHtgsWGWJ/4QoJngZ7kEgoq3IZhsDGao/KzUNHKBxGNBsQ4tN
E1eN6P7/stvMfvrAFaQfOiQM5kYBzR85Lycuvx7GpQdbK/f0xlKJ9yX4pbtz5coe
ZSWszj2D+FytYr+BpozuJ0/T3FMSQBnUn6P94EtuvI4hwzL+ZVZashJRZ39lJKdz
kZodKZkQoktgF++jeip931HxcdNNJfbeGK1Z/Wey6XisHfKq3I/MYYLWf3yjNKMg
sR2ICHQJ3tGdGnwHNfKGpF+Zlla9DLYwB7Q3XxXFGtsU38Foutwq6eEhfHhSVAvr
pxhRvgTnmgwDK9vKaj0IYydroWiytLxA9tHxu08+1FApU5QKLfY4ikBYAAUevy82
xZP+zDcF2oG9FwwVqQE21NZn+ETOj4ZByOl3iuMmIJKU5GdzJFwE5C60mVTKU8/I
KLwRGs4pIyM5gVPRECPl0GSrgLlyOUaRo4XmlgDQ8g8=
`protect END_PROTECTED
