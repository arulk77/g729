`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xp0w3VmwgyXMje8RzUirwLxZffx8iruofLGG41nr3v5Oia0tRm4m3FBtp0VEEHZJ
CHGbFyk+K2AURPU0rbHI4Q4NnQb/JDm7oJBG9PlDPXDhP0XuE7DJET5fEgeWAhmX
eWzsIDwSQtSCJ3LSXoILUZkHnMWlbbjxMJucepAvuZSSQifU1H6qW/8exx2KWXfH
9NoYuwNSa+e6uqufy675tsUDdX13uK/4ye8XPQH2hSsdifff0HT0C9oIglPJGJB1
A0PTYcnrOL4NZxQXv1sj40hBdowus/E+LztpVdfFcxH9zb8Uv5W7WyL67W+yVQ6R
t0WiOh0dL969JG0dvR3Hdh+o13omcnO7W4TW1sQcEd6EgIDDt4kOiwg1tpVNlrOL
`protect END_PROTECTED
