`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFtDQn53NZ67HdoLUs6Vo45sV5mtl9lahX9wddf+Qe8k
O2r2BQ5sgpuD4iH9Uo4qNZl4Kkz0fZQQOxCdcynfkjAtRLCbatjWlIp0XzmRIgbb
e9scLw7uksnaB1Xk2BFCLkiT7ARs+4Zk2OB/ezVw8vVJnkVu6On6KJCcUZ+xlmfO
nAbAhpNpNGTssfNMK7haEA==
`protect END_PROTECTED
