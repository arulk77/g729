`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqp4CXiBV5+kIwFXzU7TWYAXLWPEL/GH+ru/knmFIDyfL
jLvmqUuq9khm82P0tfFowk2aubWkRBSSmDh2twPuUSv/NyLMyXnsD/ZzXTRGmDIb
l7pv/tgmo1zW1jQdSv/0PGgED24iOhJl5WDXYQPwuMP5AyYlS2wxPc4UsmJnEJYA
UIkpvKtGqNV7VNOv+yzlcu1zO6sNVyqGiQzh7rTEssUEe+vzem1CxhG/Xug9KoMi
lZd3lBvRKH7fjWVDEgVyTllSpv1jFKFud2SXFsq6HzSD3VD9vF+7HViA52yPe8MU
+eMbOC8Bbol0+4MZJPpakAqNgV3L/ovBzSEkl6kRKKezcH0MuNlsRJo1981J3XyD
V9KxPR0cLP8+YoTDs7AtCm42jIrrc0syISu5TNgUqp4=
`protect END_PROTECTED
