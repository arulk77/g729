`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49e61IGf0kXtxPg6Tte/NFn8EuYIn1OwboXDvkirJ/J8
VaLyv0PsTAwJaO5PB9vyjQvNsh5wVUWRxKRELj0Igbt3q1IiFjiAka4hbqhs3Z3d
zmIRD1PS4+epuGjySoSChriEnIQ8AHloe74AMwQM1Qh8VHUa4rihgDXbNw21/1ZF
ZXpigiXQNyGms6ycj2CgjHH8wVLf7+KI05ZL/kjDwjy56TlLJ5D5xb32zNTDgt4B
ID4ZNwVJavPfLCt4glJoexQkGsnwPjNPsge38HAdJeh1ikgydGkuqiZrf4UFIxz2
lT0FboKZ+2AC/opfPsaBEw==
`protect END_PROTECTED
