`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
A1rKw93qdTVLmv96+2D1dMyr6frt0uqpnaygSGGBURmdfGi5/OriCTzFVn4nlke9
x4yURfsDVIdeORWZGYPATvFuLS14XesferXOllHRQ6M7LXqzfvdpRF96RJKMy6eU
HdwU7I9Q2zMDMCrwP41F0nytF7sBhoWLKnFE1NpSI28H+aU0woNKSYRnciXjgIvE
X6OwrHHDMhG8stLeovRdxKEw7eVEI1IjN/CHNjzp/GiRjiYplMzVZPSU0AxW3CAb
2ibOCzlsvjRQ2923bEJE6b/oA9Hn3yqsKh1iHeLlHOIXCeyf0iUgDitnZr0HcCDO
urnJu32+nlxIksJLFsZPLhvPvEKYAae/rY3To/DTdfUj0x0u1yeuvRAakYXwGxKm
kMNtJOGxfZaYLDOTyj4tfwynP0rsApRIZvNMfo97ZuU=
`protect END_PROTECTED
