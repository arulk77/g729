`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
e9RP4zjcDWzr9CcRi14rV3XniCJy7p74XvoTbk4w1LoGFkSVCcI2FvuyGFUpus11
kSwvrX1WJ1hPExVgroWO5vnjZoo2vTGdjYUxWKcPCM16vSDhqI+FvHTnxas/p54I
2VpR1PeaPdjYw35TcQyUktdpsfjeAA/KialbvHXy9zIyFWzzbhKMDPX3SLROqbGB
`protect END_PROTECTED
