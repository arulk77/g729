`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40Z7WicWsJ0cvouKPch/zTKSJLCJwR61KOlFn305c78D
Q6mm+JiYFXfcfEr4Bifi22PQZUHxhV4UUt/FKr+OHwpiRbLZ+1sC8593jZOjpZM+
bNjg6Ya1skgiovAnW1+fy2Bw3Lpz+biEm7oeWT4V3BnzlV7uxWCiXel3CTX+5hOL
V1KYDu/m1iINKNrVzGavXqUBdWHyz6bLjxVOJ8GIA0ExBWyrxyAFuJ1Goz5QUzWC
KLXIB4aOaXfkWzJO81Z1CJ4wTj8Zqc6VFx6/typM2kSZal5wE8HfdBvy/ozQLWgO
ZMF4YosfIZEG3URkLNutLYEgJeC8QWkrdilAJF17TTiTizVgllm+D+HKRzWMA6EJ
BtfeIjRbLsaH8EC40j8kZA==
`protect END_PROTECTED
