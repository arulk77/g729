`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
b+2AGI9b6HT4k5oWC90G9r2KkcKi6keVc2ibZFD95f5laX28Mz+il2Yx90PsBTfY
K5b9F9GwsekL8bnYzumONip5ZIuWP2ZmGyMerQsYDdDQzNIetR3GIDdTn/Suae2P
0sfFTU98qBnbwxGPWXenodPbkPxXltOg168lDy7sTPQ4dZ02Fb8Hqgg7va9OIFmB
LiKSxfT2Sl0JwJjviSYzMokdEM3pnMOVAuLrctmXdBnoCAICJ7mBSodHi4Q+EelW
Hhs4NmQPm7D0vaIwXgwFwZX01691UZ3hw3UYxrLefYS6DIYGkuo2iChR4DkHyysm
UvWeyENgBnQgB971SH9JRnnKHTyKgH7BroZE9w/6DnBtLnSkJ+HTTHpCPfeQTHwd
sNGv1TL+LLXgAl2qt90iRrOhKylVC6h2+I7OLepfPKf6yNQmOcEDscawarWYMIgm
uFyJCZxxBF3qMAchd6T1NYGndWePp4N1Tw2OrrcmnmJfL8vPTfscyYNGWl+BcBZF
L9ShwPYe54mhin1HEXPsz5J/ruvw9CvVjpWKg5DRSaEfwcSWdsnmXrCyFs/eh3ce
jhPVBZA7ZwLXWBHDyvPifhFDYB7jJBogTQYiRu/cvBYyepKFlKLVQnJPPOCFfxHe
OmpK6D9bVjExmjWXVDHuvnC77AUDN+kho3zZZ3joxfLLg/Zh+jz4zqTqZxR1RfBk
85EKtxdTtBZXn065Ut8bPnkCj4J9fTXE1CFC3cFzm80Jy4pJkS/oK1p73hZ7WHuJ
gsirG6NqgRdIDhFb9abJp1t7W4rmgMZS5go+zV3LJyLQI2HlxAjqA4xeuVYvvKQ+
AoBvOPM0eEYH4EvsGtuqnzPVlTvf56Nw0ZkkkEVIGQ+hwarY86pOS3KmA4K3dpG0
M7PkI87j7W7QC52rM7j0JJBtS0Hy7EcwVP9XUlA5t8133gjOmFLWNMxlsvDy7m9Z
c+fRInLUWPRrrw1+kltNj8wRnsZNF/BjlirWfReJbRC3EhTeYDuv0r4KtIRzQMOs
P7so7yMd7sr9q2bVJBPdPXin2iuyhLR5FgbWGLNC3jiAdyISTymRBfTXf+UK9T01
+SXe7ZR15hRUSZzkeYg7Y3jL2Qx2eQSTRD3PvA8RH+AdMEnehWN1dnuVgK5TI0vz
dasFApcDVFnPNMTSliShsxG9kyrAjxiAeB5EHMnVHxzeMeQcaarWUMDi8hCgxuHb
tW1shLihkCNujb8c1u3gjq3owHlOT18WjuFbLIDvy/EgVRo9vgBv2yMKQtHCZk9u
E1mlagWauOiCwfOtd+RHWv1VnLSbSlTaeL8G02SJa1qAsEe9+9/D3WnQPvTyISne
uMolhCDVqRBlYLx5Zyd+FRPRJHUUsvLG6kCzp55yiFGTJ9bED4Q0FfA9DaHKpPJo
enKT8mPiPSSq+sCExiMbF8umz4zXLoPRFhvyJX1lAvGow4q3KdWzwELVtLSRaYyk
5mFV+G0iA8iBG6Gyp6fK0CdL6rIz2Gdvjizbd2CJHghYocMtlA/WjoiS67Ljji3A
g3+LtBM7CK9FdvTsIChYCEYFoHtYtXkR5ToUciRSgV4elFKy9YaGOQlGGqJbxPcV
d3dZc5MVteB8HMHNFHUpew9RJxc0W40rgKZ7nCQmfVMwbqvpe9wkWqxpxKy0PDT9
Svnls5AlZUae3AIV0vbFctD1ZURm70h7MM6jtftX0ChCO5Xe5hDMx/x7XZTH6t20
gb1xRmM5d8YUCGqeav3zLHtRSEZ4oCY0T4NPdSol58/HlnrhWRJhzMfUPx8q0YzF
e3Docc6n1G+kJQX1MGdI1w2G9sI8lu4cvkZNWeFbPNVMKU7EMB4lSQZtUfCPZ7Gr
COSNpVr94lOo4RZS7jaGeNHpH+RTRhyfJltgyzXVi+1hKwlscAUKyJUiAwyyXGtZ
zjfXAJ6mMKKxaZaoC8i98qP8P2K2wBuMkFGZS5af+JIFwbi6nrfwRAPT0MsVfHs3
24i1Vr0TD9rnlDJ6Mq8MPo52froU4VqL+Ayin8ypf6IeBN+joXX0+w1mV9Wh3A5p
SjjRhJWFG6P8qozP4zsIiXFmyVvWqsgGuAJOlGle/cVwALHBSIuEDxuggV7QcE77
ki2agWxg0LSU5ZxeXtg001SzA+EmfdkwCOqZLPi4tUbWGTwUjGc8XSgCzYEm5xBn
uQNIzk+5ReSVpr6gimUt+Z2uAAC0d7zdbgOEllifLUgoisnNCQr1GB7cYsSDvLE8
mIBOcuvqovepRge/LU55DY3HMUY8YDE1JWhA5HI91DJ/NCx8TAly7hg8dqIsGfI1
OhK4+EQOQJBsvQqdXThUugL9Uy14yZwQ2DCEBWF26Uq7e3SYpyikJCwtWziPsE8b
iCdvHObmGGa+fkWU+TkEYQCx9uaydCm7T/JFmBM8h5x0jjaPTusQC9785TAcHZLd
rFV9HfKG0eLOuY9oRell++xoSStvMC0wF+TkEIknduwpfJotc0YEjRcP3j1NNp8Y
x1FyKXSry3XXcODzndygvsv8WI5GHE4rFoOYR6UINCTMl/JiP2s9av1TXsrbUYS4
fr1QYvHizi3OsRzapyXWhEhmyTDKFdzDKgNiHNnkO5m/AVbFFtdCAII3WPBnxiJ/
FwJIa84AkTUF0YF1TiYgYVviugM2A0WYcwyw4RK8eIMbS/i130gRF4MDPjIGBTkR
LwNNBF7YSwRQw7SprFLDPVJur4hGbn0Qu6rOGBVMHCOAYFAEr1VG+3spjIcPJKEF
t2d+dQmac5EI8b62Gk4tALVf5TcAA10UE8YWLjbCZ4s9I1G3Y/Td4FwEUMCvOixr
PlgKIESthidJ1SGlAuMnJD3NwHhqp9HzxrxIzIeWMFTsMVyjYDozMj5vGOO2o5V/
/en4N9sr/R9MsN1F9AeLohzZ0+RDViq09+wjx7HxzeUQMiSwAf3Hscs2n180qIPz
DgC6kzpva+hHD+OHct/ZsQ1BiTDZp65EN4SclYFHfVnW7vMaiMoHsECcxIDW7JUx
Kk9tegV5YpFH0s3XyaF7ugSGGvQk55kdx5IKPp3whzjKCkT7QdIrZa/tvBpwRG6g
/dov9HkUDt4O6lAGz14wdIY90ENsJfAc4Rj+pOzIrTt7fqEq0/hKysPnx+HNVnPC
Aq8F3+O3jno3Xb/4nFcjFDNTHU5C19DuthjUjbqUnurV1lpHKhvCBYIu8EOxN31s
tpU1bKUdWq7uDdwfZ3MHG3WzEJO/1vrRTCfgX/1RTibbquvXyjXR+/2IEVnw9qgZ
Phltmp5nQybYi7PPj/1kS8sAo3ZZHC7iZc4gGLNfe/3Qq6g0OVM/G5Ha2eTqYz/o
rTTCi2diQ/eeDsiSmpfA1hR9C/0AJwvjXcRyG8ms88Ae3Ft7mjhlGs2+lhF3lw4g
y8iPIKfEQVesvDsjuhkbkNoRA6snIDx0hLAz9CJhFzj6ZVZpVaCsRa4u04GUT2A4
6qKt9BzINizaGu6fboHt9B36GJikDi5n0RwVN3kAs8MldDYbtCgteVeeFejc7Fau
9mUNW3vOMEI3JyJVl3OzY4s2fswn4+zFSjh0L8oZDHu9D5G7LPS0YCFmgYV/N70B
0tmPbtus2Nrr2yz9AI9Bst6IZq94W1POw8iRe66sJpIgdf0Zplm1WyECnmGO9UZn
jGvbRx8AqiXoGGy7N/eGdES40qFJEb4t5b69JJ0V4s4LEsWMDaGT/nVhXhKyvWuS
fEST9zsADfZIc0IFlE+6gb6luxNtxqhvqRf7ILQgzgssQ0YWWw3NbJnbPk5xd8wC
YEiaWkZsv0daGFItngLGA4XVtPnJ/VQD4fd+AWjTZEF/93gZ88l0PMigfAIysTVS
xdXZgovdajaC3dDijpjHsDqYBEdylvWZorpLcppNSCCu0uQ6clPFfc7USOZOSOAn
ipiKfyXjVsVyxRZ8jQTJ+L2pF0RTPriOoxmU86em+YAhknVZmxQ9YUnN++vWcU3O
Bv6Q3JPjybFJhRdeeh2VDG786xfI6pZRgolZTnsJ2MCn6rOtZgiBWPTAlk1DP6G+
iXDt1SzCSxFQ485DCmf4YzkralEEfMnIZFnVDHFhSJ41vmUa2hx4K2QibEyhS3T+
6iXwZoyNd12LyDaTN/A9mFYU2DpkMqCM+K5y8ZTgGfVrHtP21Fza8/m4Wrs3+Lrb
AsBg93Q1RN6gHdsLNgqntLWvBQP7Lhsrq63WCzb2QHxx9b9DpWo1sNK8kDjhL9xl
jiGAbYZL9G+O3TT3nriGmjYPq2v3Th2LJ+DkbRnl96Z5g/cAwRL1bOHOJyOY0UcD
GfO6xcT8Mv1UoFR+yJB9Ctuix8p+Cmj7abkOI7AVVqm/yvFX60LWj2GzJ4o98gsY
MxEzrUiwItxHdvxQCdj4rQVjNh3sHxDRrRQbUhwMs1pgAWh74iyoK9XiiBFTJQYd
pSSNyhitW9bsDQCamO7Vb655TMwhZNkaTPHHyvlceQIjj7IoWOBVxO0wQdOxY2mg
RPqslBrXDZ0SDRzfU2FvXLQhH/mT7BBiWq+M/zXHG50jlDPl9sZZqttj2rqwkxAV
lxt6ui6VxO4kJw1D7lQhe7H3BSF2gdHpuhxaQaqg0RddMQulP0+U0HSYz8pKOt1S
8+A6NP6I/YAmr/Z27+BM3nwTzRMZiqnKLQNyjf1PM2O5eLXpNztN586QZc40HZ/I
pJanI/BjUl8d/DGAvOPt2bHtdHSHI/l1D06PmhCCZzPgHHBSzajUmH39/w1iqJsS
uNeQG+8CYk84OPw/hH/WDWogs8XU21hdCy689lwfQx9dq2h6bc6cCWvSGOfm/0d2
wAUmCbLtKoRQ09+FYuOAzuxN/RdP2eVEhCebWPDslUZCwp2Ye0JnwlbBd4WxBX2N
7c54BbBQXr0hhBNBX4gcfXu0xNsxWcSNOpWYza7IYhJ6Q870DFF83pWaM1iMBL9+
OyeirX9DaYTa4UPjM9/3KsGIERVu8DXAIp7yXraNz7u7ECrCQPWOjpiJeRrlftNo
xAZULCH9PUcx/0nzHr3yMm9rrwPjDVzVrUcKobpu/evt9uiCk2vXy41PAdvnM/E7
bFziRjzm/L9whls/YYN2cGqLK29j4pvdDTyaNRVcynBAwqrf3gQsMlbdCmt/4bbK
QMi4BZgKPV+kMSr7471IwazrX3lBQxOls28OCOqtNxNNA0/hmOCFlSaQ/IP7SE0T
LOv5dghO+66bVur7P8+ucRrHnCWndrGg8x/xR7A/10lgn54lF72HZ0gFgREQohQ9
FXueguT+e6ADZKn9hWEOET+1sHOXIBSU0NfrxpDfdob3eJempz8MDljIfpKz1eA9
U5A+AOQjVkHRTTw+hW2L7myddV253hJJWoU6hzn59jSyS7g5C8f3KA2GH2hXuj1C
HYrxaNo8qUMalDX9w+57r5+CyGycaIpTePzVuO5TOLIQKLYpthkjCOf6YUsvdaoL
Fw5HDrZz2/g+noRN4quf9N+7EgTPqeYgudZFCf9uWSkQFx/51wUO9art1V08Lt94
Nq/kdh9sPCvXPqLKsGXpWql1ZIseARWBGFD7qkATIzFQ/kQZjIBh0vfuu6sooWBG
cBCnQsI6V0OZ/yXCrRoYi68qOCxyVxytvIgqB8dQupB+w+6f4t4yzJbRKFXlJ/zt
Pl1pGvRYnkuBbWtNbdD2vMJYrklxXYL9sRn3nmMcCUhr4WrKHD+0xbUvQ4sp97Ft
zo6l28WeFG7WtCulkv9/fXJGIqGY5duFzHPeyYu88nWy6E2dbuXg7PTGN6b3Oa9K
GL1osrBiMqeAqihjHTwD6YqLhlfoog+NXeUQEfqr4nZB84k0Wycs7Qo+LroIBUSc
gvQnkcNqoYtRMKQfMxospjN0Dp46oplhDqAfs+jetp6L9UGDVLknzVsdgCV0Bn5L
vIKu9U6yI4Z77XZ51uI+6PMyTYLLX8SrEQOpFizRMqhOW0wKTjZqiup3jzEllOs6
7ZEsuyCjeMzwc2ULfEn6irCeNgNafg266pTYALC8jDxPTCv6bVSl2mDMRQPWRQGn
u7Va2l7CqnWeCaupc2FHhGoTFJH01E6aI75AoP5kHdhqFxxreyFIuJqcyBpInk3K
Z5GHYDD/rtGKL014G5ETq+Kf19XaMsGJR8P7VpN03bibvAraq2hwuebPgdVJ/qId
RDixKCQllZB4ChEw6eYX9//S72ewJDHxv9IKDN9G0jYD5Wab3Bmjdbr5oyDnLUY5
3dlkaz8jZOATdjwsCvyzPxdACwW3At2skg7QXXWEQIogX3sPpBIqBapArP17CJsU
Q0rAQeyz5izGSZY6XCiNfcn6iHg4UD3bSNi4aALCURjaDWmwgOKSRr+3fnICYd+K
Jy6GdyH2y3SXm1q9QemdSNHOXuD3au8L22vZbE9HnDVYce4IZ2R2dz3nDxwguQ9m
nD4fVXkn2+LfNcQEVyP5Q5jKVH1x39393vZwArpTajjEtWSwRp9i2zjY5AJ18M1s
7RgdxT7EXdrMGdroTaHG9aTNZ+jw8xtmwJW6nTPcosONuGUcVdoSVbsyM36Tc9IC
xvDloaimieTHLpOPtC4UJhK8n1lPRLYUtOyJjXajEqNC/XEM3toPS9Hq5hDm+AjU
`protect END_PROTECTED
