`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF4haDZPIYwIEKqIVU0tTEvp0uzOjap7L3YzNPuSY4Xq
b2y+XGSmTb//887vXdcmSZu+MnYEsoFF5L9vna3JW9YymORhO7EzffvfKTpWUaXS
3K5fvEnvvzoC8T6KMyyUQjBh6Y4IAijGGaHgJXvOj/pvm4wl6ZILKNOOvEzMSGHN
7dRxGHuntvAaQe/Vdj7QHQ==
`protect END_PROTECTED
