`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAeGoyA7b5+Zl4IqVvL8KMHyYl9I0l9G57hUZpDFjNlxB
TyUJYWL2Gul4j0b238MyfE1SjhoTQEvFGUJHCnbJpfX4PL0ii4iYy9btXS/ks8Py
ug/nQs4bLQdNkSHpuOY28MW0xMUJgC5wRgTKp+5GcyQbmBPxNus3pVdMFNvXoirz
dsuTLr6ousdr2epvr8po2Vk8Qmnnnf0Q7HguH1rSl2w2HwQk0VeE3pnPUnafcgDO
t2ki62pettnkdcyCNAmGp6kbyFaDXuPBXyeVHZusDNhVOhAiHpSJeAiqo3zONQJD
Id9vPP1zRJoKjoJV4QB5Jz773iU6EkmRrwPn8k5Ltvg1vhjA3310inguyVbk+Nm8
UXUfFQGZrOFA1RBaNUL+AI4ehdMCvyjY/LSW1d/+xqEixNwll3xVLfk75Qaqr1YU
nqPaIFL4IFkpQF+6yDQf80n85OA8yFhePMSOfcPyGEkeiHVDjN+plermJJqiQ5V8
bfNkkYo1oydamLS2XBBb+1rGwQYqIbsGzSTbRqyt0j8ETohbu3ZUalOmvYUdpNVd
YWRYPwABg+53gtA2QpODV/+U71Pf/5KUKkiRaKU31M8psR/JdIgi6KwNqS9skqri
IkzdEv9JWFLdFJVkT+zsppzp4/+6mCMhTjoxdbSSnlecfDyLjQBQOwJiocd/byi0
3Af34V4RwLvr24T9kwva1x+/u3Sbm8w+6FHpH0kMa7dbPOnYhMw0iLRBHQXRP67x
vlHaLmIRdXTpo5IJidoKneErqqt/lIGIZs01hJrvKaVOBJfFyBc8MNjOcpGgz/sU
Vy+lfRA3c32OTFHrHrohAF19qXthV93wYpNmd9gimkO4TU1Q+DpBi0Dx9ZSQZdoa
f5a3qzK+xm543jXvrD3WXzB9Sls+SZycki5gUhaEBS4etjCU6gVCLjh9awn6n6n7
Vpo2DTyrFk2XpwQI9UKZVZebCQgLQF6cHu9p4CRv1E+5Atrfv1n18JMwGi2n8uQs
YJaUkBLhopCGTkEw35t5QkijXSBV8uXW9Rl9HkApJ3ZQg7ZEYcifblqYyn9VtTpd
iCGYTOTpEN7Uiuhx3vt/lk3DCgzv7aiSLZccQGB7xUob+njiAmWehLRm2pbbMRUF
jRzV/SdvRMXJnkNlMYFZbuPuyUevRYth0OdkXwWtbgPd+S2czkZQFS3bqZdwe8MD
OEjyn1FSKtOvEd0LOZwGChDjWGCFOI9a+eNudtUIsDNbQdoku9VRZ6XWlT/qL6Ii
q28Bql8pYVq5YyVYJuzvxGsWR7ckhBbWNGROfrlOVtx/2v81ds//T5TsJAoq/tML
UPnmbvpuX1ZzLsYoC1K6weLNOaDhpY2W5BbFmmWxRkyRZti3jDB7D5jguORerpuD
XXC/gjFDnxbOPh6n2QtE2bz7uq12T5xq4RCG+5hCANtY/yn9tyys59yEu56Qc+dg
TnuoOqKLKsKCY8F/+BFKDhFuh137e+R+ozY+eKk9aDY1KO5P2WUGGFINNWIFU3uf
uVJXraBasBnYBNyNxWscaIbkEx/1x7cnoadazrM+kE2vizLXPYr2Zj/yZ/8vXpqH
ys2szWLCeoJzgF0YCXgcVl62PCpmxBm0gAW0yhFmnPXLHEu01u/00RANcIHfVB6v
4jImuD4NBTSEBQajS8nGrWVftrM+LEj9/KkNHpFIE5lm7BHrMeM5g8ljTyf+j/T+
8yfQiJzoWhJFDnhuE58QWPuO2a3wN6DYJ75MsbWKy4W/u3s5e6MpNQzTLao7KMuy
eKGdc8PBRJAdAzlsvkSB5Iz04iGbonAs13ZbMHUv0ftq3uHVddPOXlLjkh32r+Rt
DkG4XcDXNPZ7oVOtd7nMSBnLqnxFkGHrEJJcltenhju/wupV5Gv6RBRDw2Qto/dq
ACBhtmU5xQbye4S/0cPY3kF6uTJWTzUereHXXbvtpmDvP6VVGAe9FYEiDm2KduTU
NIPTdRfgDtfIyiuHSgoBqitcNg8trCqwTDC6C4dLwCOyTVLV3r97e1E4RitvQ4ZX
s/RjAQSu4DJ1T4UAA2SpepQWzWYmqoun1qq3y2K5EBLybxCrWRVcp215drBaCxiO
eHnOCIi7pksBWeFad0LI3lfCYdtivSvXxgcNsvc4Efw1Y+NflVHDw2axCkZcKRMj
hxwtoWjcy/PlGnAWV8pUbh2Tnc5bCZCtTclA4WFjY19WQ6S2EkkdbYLsp/nORamS
veVnkU5hpYGOSmvHPbBL9xuuXbV/IqxMl4ltjDb6Sf5oIiIaxJ5AJxFBgOlhcIiq
EmL+iRGFot/EEGQ8tCkKZEWMEtZZnpQyw48XPjNupOISKMCiUe7OuuKDbshWwzdL
FkOcnqG4/MZ/V8cytsbCiLgGqYXfycF/tQ7eeZPW83d71oTt9z5T8wD/o749OvFq
PAIma8b75lVFtvBSyX60Vh4Zn/ZZxM8jgKzXCDsxw+FFf+8JlOxYinXEtm8s7Kfu
6eIoGF781CKZySPwsOqsQuEXMbTrFdBK0XXtvQprwPEi10RXIUWwbBxpb2CZSz5L
U8ygEhU5hsxnCTIvZdyEpI0gwsr8eHMU3rsnvuaKAoePBhwVmpdOCqgbBXiJRWUt
WA4Bau9xzhEwqED4CGLdAPWvgOPEkEgx6uo14cqdcXkphau230bOp0TPbTblwjcQ
xKxgF2es+fs5B5WOWQeud9phTtMTg7iBK4qwMqfmua1SyNgZtjIZNc5PmpM+3NIk
1u2EQpj26tvTM6p791F2iuktaq2vWpGD+dF4VPHM3Dui8i6OHKf5h1TS5YD+hPBz
K2wRKFBSBc4U6I1tLQ0V+c+AKmvMZEYBLkNnE3rVH9xl6MScTviNHxLbujiaxVzx
dFF/vLqeUYpoMi7e+ZV2YMfVHBo47NKtP7+PTrL5pM8Fwu2ajVd7qK2H5Opzrd28
M7RXmX+m9xt74EkrtkvRQJp8djkqf3mrfYOgZMv1o1K7DFHX/arwAb886feheaAG
L70lE698AuvGmIHstb2ZAQSSd1WFYYOWqTxQQ+gneSb3KEwOdODnEYSiTlla3lFX
oMopxyaI3UQD09qD/22i2knT6NLauoUF4TW6rD9Oqwc0qOHm/DvVkHKqH8Q9DY7U
evcXvWUfW/T2dmDUjL4aE+bk181t0LHSc6sw8EXXNf4dNvRDiyb81AuDN83jH6SY
k6T2S07ewi1F5g4JfN8EghAZ2oY3bHFnGB4UYXQNSkjoZ97DMjgstHB4TaNhlstg
C10qFGgmrro9OOkMwclGN0ZCx4v2rEpvs5PvGrIrNktBIBAVZOcu/rJ/SYUF1lXf
srkmTvSUZ9TwSdKPzEZat29aRdxD5206Obkv2MsZ4v74pngNkGVbIVIFarqT1I/+
WRb7RhadUPeueLsEvyy1wVOgWoNsZnLUfrLyNbP3+b4KYewussWC+slstLg0JRjC
R5EkqPsSjsjtgT/F/fqbdqPSlYFM33chbiGpAWXH6bp73j0YHccvDbg3PjnUIaAM
xcOwBYBWx6UFh7PhxzyDjuZ35PmbDeoF0YfbJmbc9kaYAoZ9azN1PadPP3Amd7KJ
XsEtQ44IomPDqogmOPvpM8Jp8KevyQvneadG5eE2PwpdGt2AnGfDMr5IIz691OzR
9k1m0tlIwQknX7wlisjl5C04NAh2AopixBBgs3oVCBTQBMzV8WnkGS/Jn7WIfIUD
qGZTIvhwAO/MHH6Go1KFo0dYOqiLEnNtLnvCTZFruuGF06+fPG0eHlds159YA1VT
fhhUULeRD4PHjvj0kqLx0TCDNwhKSNx2KP8hgE49gAOpD1uS/RsU2NwuXyseus4X
XSFVsqs96E/G12vHhR4Dg+/Lg2kSQ9WROwqDYNce6qBIQ1JOe9DPwy9yrwu5GZyo
PBG6Gd/iS11/x7ELX2WWarzaHJU6F/3cw4zCsRyH0Q0Na+iKZ4c6ZWwog5DTgU2Y
K2YeH63UBCd6jlfIc3HSpSPj2c8b+YtDjupSG4H3aQzr2u+Z86Ndz8yg7mwqCvpj
afb28x1pWfwAdmSJurd2tXlGFLKN5AL+8mypvD6CxjVjs/vgaiDl34lAL5qQIVj/
5vH+NussfU1j8dTuRirxKTvgAMnrEbFBJnwLV1zhrhrISBcm81KNMf1iPsR7Z+rX
uJar7IF5+RNo2woRlryIrqQ4rsleKwKa6Ce4LQfy9XUFJn3+gCVo6VXkAkn4ZXPS
5x6TRUqnp6VutGME1NKauVxciPImx2LHqYVr5fCFEBaw4PBLbkduSogkkwp8DsZI
llqbCq/XeCiSrnem5qSdSF66YMVMA03WcAos7Jan6es7BY9DLYU6S6cAmpH5WLzw
snOmVKoadY0+YX5Df4V1i1VlfsPVW8A9GJi+JBHbA+WhQXYBm2YiRehf2pzgJ8IJ
u0YDhxkAFyEChpUsA6LlAHwxj8wpFsnDrTg4nqJOEmg2pI/8Nze5tuaz1o35nv9h
kdCykvFLA8hsLiqNyfpHAbkaFEqXBhpyb4RUQfRmnElMd5xDITnS42ShxRYMLIK4
6mfoFgkDDXDrCi37H9XsRotqagxQuIKLK8oL1HKsV3wjd9JOCfSmYu2G1BGTpUKD
504YLIk30oBHxyYhj8iNSonPygG+H7bu6HWqjDn3lr+UelXtCFKWfIkFJBNShCWc
6oWVSvC0ru/fTepxfQw0yWNJWEZ5XNzSgSPvdNvQgBLnWhO6fhKfP94kE63lpo2C
P4hTsjYN2ODLWQg5Zpwk4YBTNCKg4VdO8KAl6MvvB/OXkKZKOjCMVD6q4pWHgYoY
uWi9qCrEGrXWcNfTPmbO78dQMDbzjJfs82gjN+FkdTkIVEs9mp3uiMxlauvKeG5I
sX8HLIZgvK6Xqe3k/uTKqz/S0OZSOuoE6xPyEp9c9bbV2Oh6JxXo3DAGVHA1iTzO
8O5EnE4TjM3YjbCx8+7FHd14OT2YKq/bAtMSK/1w7A70oTVgTkGOu5y9/s7m1oV4
iVKOx6jZ4HVef2xzXGcYh/aZ9s7KrN16FALUixG+m0h1ns6GP3REWpLhfnB7cPzg
5Ll0obHLFi/ygkxRRmlO3IWk01CW50ZVfmMd6HoocN4SetYJlkboe2XsDE3A6fKX
xJh6mSJWNL1ffROb7Rl5o7J5stRfeG+wMSNqJVlFO1KIMHuBcxqemXYL5GqHQVc0
e+uupf62agaCWPZQ9BU2c0HK4BtDDwAKnwYA3x8dS5hsW6Mkmh60X/kBisQDSsmC
2ClkamAr7pMFDVrQZpAO/Gx3WAl3bC0n5zX5BXYiI7kfWdoAwM9Ah6OqatSm09gH
GOBfNLbX7Urk1uX0DpclVvQB4UOLIBLUdIE+E2jPCRU9rTmsIt8KcFmcDeXN3D6H
v3uF/+LLE1MorijWF+sxS7iblUTWB0AXvz1U4wwDou8np08lPiRkOiQlea6eyOUg
JD0vYDtSbnsUKQyAUv52UxoruNqi00KDOa6mbS9b/fPOYUHjzyexfPyV8qJWn5Xu
0VpRtDV99duwJkxrxLTZkJ1p9IQ0gLYx0n8N/HLF58KgRGveb0L1P6dW2fAN2bbP
bwwfs4n7sCmt8Kf2IGu2QYGylqC7NgJYlzbfTjgMEHmgM7mkfG6kKG0KVagvDmCL
L7cyv4qh09AfwiGYu9o0smYm/d9uZKbj4BlcBW3iq3JgkTOhG1MDJq8Y/Cjodvtc
XVNnhEiroYTSHKyVvpu1hbIMPz+2RqUKA2e4ku+/K3m15pGo4rmmiPDcNukVk+Su
LfJL4zHcvtOnQOBPJRnvD/+mXkruF4Vs7utlFAWcrGj5vtUVaK3PghgMbg6edYQG
/V+wMcbzI41ymGTUP1byuHa/j+igtABb67g7CRyK7WeSWaunMLb2xA/goIgprbVl
70RyPYq8/2+SQQWvAprsfq2fv75nNHA6bYYsCmLQ2nE8N9JnhwXYcV82JIDClwbQ
j0xt8oDQEmbs1CfthCzBJirJdJ6sqX4eFM9dyWIYWV4wwpXur5MgfdXVhldVwM38
tphZiPXc97T0Nx595xOoR3Kp1vXo6t0Ibvt8QC8VV0fkyhrso5dbAK+qB+IN2Czc
5aO33S8ZQNBEE717wKlH2MZU7Uju9jmimCjPNuzAwiV99/3k8GoDiur6EXspX1YI
o2SmlqWMu4ssZ4oCjIHWKPLeANMKtMizxem36+g980qwJL+6Q5FehSEPCNCEyIja
Dychwa7L4n5S985NCjNNCT4vhxaBoGiigeWZFST6sCiPiWtoikJLMZ/z48p+f33V
Z5itYMpaCNl4Lm6MY794exiorsrIVNxETMjnSSh85LaK9eW8sepcHeI8qCciUF8a
HyvamG45Iuji/yb2UEfweTRfvwUwQrjGuW5Eidz7bBLwO1zbc6BpL6tI7ugPV8Vg
8VYrRxwLTSfjd31JOfk/R9c1zfyBiRZ19BKkagxcIYKNJurLFIP/aY2Uytb43jsf
MXp8mV0wINxlJoITQvjXy/ZuHEay8aM31V1aymHgx8wgz35bJ5VDQBuMeG7vrkP9
mkevE8SzHPsclihCtbv5EPFNeEYgBShHBIHwIvOSxZxeanhl4zCy7VY+IF40xPGx
GeduV3HG2lfdE1P7my2WuIEUTOtuud7aFmRKdqLyBYMhx0IjHsFGbJ882ospfEij
qTc/nBwdUxBkEQcWgfemZrsngQ+BjF36qjWt6bC7PY303u51nQB9J1S3wV1wQ6XU
leJSNjHQhmObspqLw6JzIDCI6kfeVU4PYFMoGDb++GeDTFh4kdqu3MQA8TXRNqVL
VeW3zWhxy/f2smINfgQijZzkTiyc+vhgj9KvVVkOh3MggTLFtXVA2CSMFPO+VXUj
5/UmFj8oFrZWI1uawEY1De335Y4ep9bWuwOZV4O7OMRiGf4pKi/Ls+hI67Q6KVwX
DPW19eB617bmA3NFlYEQPBLKAZksKjWTVbEgs1xgvY4Ka2GmteLlI83d4dD8F7DC
O9Hu6yQcBi6znGk6nHw8MkkvQCS7emWS7y4CXD7rQVI9YmZrj25UAwgbL75gxMMW
W1qPhJw3fGYTucpjjjcWaIcncBPrzTO4VE1nOW0dgxpadOFp8JQst/guBL6Dxs/8
A/mLg4L7wicqKMAskiDg32oVb2JxxnFdPuaRByFQFcQaV2yANCIIzgrfIUEjDLuG
jt95P5bV0cMzzB4Dmc8lHNa35woO6UZT6Ge70H+2E+On2zwzmmD5nIyjF3fOTgfR
mIt9L5N9E9RaL3mv3ytbqTLOEM661ktslwn5zRrknwpSKG/QDLjGdqZYMDeg1GTk
/aCzdMpWH12nTE1Dte3pVfKzQFmkQbwkdfBPKTolYuLaDxmw9W/q0jqwcDyURftj
1CoC3E+AZqBN3jMjq8gKjXhOe7Lvw6vdtZz1MTJJIxPbX2ofFi2rMKJLfZbk3Iyi
I9pk183sAe+sCoCwEIboNbqhy9C16s/iqwm8btEZ+VwDIrduI5dmGHHrTc/ZEYsE
2ig8za3AWW62KFb1YeL9CEaJ36vb+11mE9CzuqlXMXY9/7WoTRlJha90pr8vZnrR
98q5rOcmBIq7+QvUPBzoEIv3nKVlB4nJIHgfe9fdhl+OdS6MJPO69BjQf0dES4wA
xm9EXyQVwFGFtyNMcFUgQ8DnYlOslnyhmBKp7auxV1G0hJOnlEQjLzWV1tCxLsta
l2WlILJ+CYJ3v0uvHPL8lihRh0O+dZCZBGmB/55bArZrnt7yQOXhBYyX/Bqww1zR
JycNRDLUllKkpOB4ZdxT6zlggqLnmY9KIaY3TCrlROWqAsSMDbduudiieu48hmo7
h3L5Q4JeN6A1XNR3f8nDP93IVvzKT9gAbG/Umkg+THnsiRZ08whgvRkG2wSAAb4i
`protect END_PROTECTED
