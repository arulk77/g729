`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42hKeFIDFbS5qKSW9HsNdNZ4jUcxBo59vQTS/BxrMK1p
GFJIlya6AcNpmUle0BstSde9pf75KMHOLtUPgaw0VKtm+H6uM7TorEXCefTpWHdw
B5MSP7pT0C2Di7m3KGfqppeWi3Xyb3J/epkI71T7XNcTugpXIDoe0y0bzvYzVWM3
R/oW2OziRrHWu2gfrX65Pix88fXMfcC0aXp+4KtlDJ0JO50rxIdQuZqcarXS+v2j
eMGvlFm2EUXJSlmqy0YuXqIWjDPcsPaPjrn6C/yaMkeik7opw9j28tN1KRMAwGE6
J5UiF1qTr1qqIXUMWQi1rAq/0GU1p5dCGM/yxmAfZF+6OEMg2wICaKjF6cMfwLdp
StH69knm1+ojaGQ9nh66BA==
`protect END_PROTECTED
