`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGka5oHMzIKvy37zCUjrLU200OabZHdfsZhNcvnKcoTu
Oyk+gWSFJb1emZyalsENjWKg4Thgo9xCJl++ARXxgjJeKP3u7VTqrW3VLdZ2UbT4
7DVXHa2X7Xph1lvpp+ktdQ9zVmJSJpxFr58uaOvzhnd+sldOjyqQez2XcviduK3M
LnbeSf1f1pvKTl5nEyNIVt1v4GjYwDMJRyiTJLtwRHPqwiSwWMnjQ0qDbe+0i6up
`protect END_PROTECTED
