`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44rqbS6wuMSgograQvoRWtEQdEcNDjLinDtScDqpR1D7
nah38+eLOE8lR/k0PcfUVXLMP/PtyTumKJtKJcWhkq+Tb/yc+kBQC1Uclc/YR1KO
CEeRbGjvNZqhKWplfZeQUZH2RQTj2edkJdyhlnODQoj3oNgjUWCa/fbnVVSiPtzA
v+E82ixSV5TV6HWOjH7nlJa/IEM3VtIHG+xjVi5JDH+BvtgGNZvY8/Z7KIKJVyVn
i/zfCjo5m43rBqdj0nHqLHIqBOgZOu6BXPJVJ+kGPnCQuSbmzWK8Uv9si3o9ADWg
/ePNT/VxyIwoXHpM4dt29Q==
`protect END_PROTECTED
