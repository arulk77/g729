`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI39s6jrmEc5W99tBhuxRFAdk4lBkWrEipX23HzyefU2
jP+6VFjoyxGcoitP7qDah4s/RloIh/kxIfwb6+9KSTdEqdhRFOSEjpbA//vLf30G
wcqy7EncXqlJYRYJzEw1p+0xjGqRwlxq71EbbQCJOp7So2hY651Z1FcvMgPCbm2D
8eScyfjhf1iskHo5Y+NK3Vv82AHLSJ9i/DTBqaCqRNwYmOQkEXnoXnk3JeJPldo0
oH7hEzk+OuM/4zlj95+SOzGVBDXE+op68mf3XKk9SRXKRqG4v/D924tAdxsWmQxc
69NemvH31vsVHSc2GAw+CX1xnPp8NpjoCLpV3apl6C9SnW/IfqQJnftNGw4S+GJ0
Y/zcQqOV1VVQXSfJbzV0qySAxt5BbqslV2+YTziGvBVGFbOM6CJsGi5zE1vvyQUg
lnI3NPvZnHgi5nkzb7OCehaBGPvFE40Ni+NhSnkGv4BCOkLBavktN9Yh7lB9JP4a
eOmxo1/OZ7HKk9zeQQrAZuhg5duS1smOr5s0+aF2Bei97Gctn7H8AV4p7lsY2I/Y
GRPJccbC0mzIAE86NzV/+g==
`protect END_PROTECTED
