`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
cuaO9m3anogVxyMeJduFVMpq0aZZ03hra1vLtqNZtIa5+grwPpwE8o09VrqmSKx4
Pu0MRJwS3gIUNVZ5ltR0YpDW/LmJ04ueIqlvdoxCKq1W9E35ahky0uO671WSPaox
uGS+eH4R44vThiBjS9ar2739cZxtlEEcOSSUWOtGxdPrUHDhF1gXE7brAl75lV/n
9x9kQBuKRCqwrvlt6GJxBDtFyStmdKz0beuKWdmaocTciRVuvrpeIK8pK57DUuja
nsSMYL76LfohpjiAtftWfiBFXPr43yTyHlMVCtvn0W9lQDMc25Hx1OujTHChiofN
3bV4n0eSsZxZAnI3WuyjolhOlroFhzJeHAW3fFPur9UvF5o1X69/1YNnAcFQXw9I
N/HwRazrq7xEMF0kMIZp80KW96FfXVLNNpzwRUiBLLtvyEhKK9pF+UZEjhr+297n
/cxHHYAQyH4d83S3b7hOa4kHw3Uas8Vq1ctcm9g3S4JEQWL+RGe1132yUXUfmFqD
wPPNkI7wFLQuHNC6sCc4As5WG7ReUqwolSBWrXcDKiI/qDsgEiNbM+eARcV6Buo+
ydvXDRpoSLSvntuu95RQAmkGqmuT4MqZ4Yx5fZiAc8xcveKQ156Out/nbQ4wZFBA
`protect END_PROTECTED
