`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45PNb/MU4SO8ytEMU04lk7oapeBhb808MdKYqibXg03+
iRntl/cAFIsL92utlzewJ68rGTHkHqBRT2b8jiZu/4A3/AOPZi9L+Wtqppr5eDNQ
Izgg+p897XK5MDoRC6r/nbmH5vZo89y+0pmJBBuDLuNLeVlI1KS0C5PcWJztIneI
liEiRwbq6nKIGc8wM8jxaGw77axhWVZaDvVLZOuZ8uOH0aYOLxZpp/b7ll0QPF3W
LJ1WdcMKpjmZmOtCSgty2Pwy+4mRgezLUxyfptgDsdQ/6HSM22gXdi8T21Cm0xAo
WiAYK7R8MEkS4GE6eQ+oLH+HN5QNFO+c543xm2LmqrXNBFjy6LHYhmNzrH5Zfdzb
MPA4QzlT0+rpChfFApPx7n9u7rJUivIwA2ZzPMjxGSE9ki++E74U4/pZadaNX//r
E+u2XzZEqk8CpTAT49PnxQ==
`protect END_PROTECTED
