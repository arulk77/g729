`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kgCJi4aYnprR9pYCLrbCRuFog99rvOJX0ymKLUnb3owRgcPxbGGxHYBeO0yRqYTo
HC4C552kOkUjtcLX1uAVMS9ozByZodVsoXZS4lHMiWNqMAy4pBRQgazJZ3wrnTn2
fv74lAVkdRJpUXZ1lgSVFBE+BWhJZOr/On1MMmtB0fodTs2g2hblV+B7yI1eUR5g
eqt88Ct9JZzP+VFqInZRK4MhYSx84DV+S3mEWxkwFN9oKE0Js6GmUtNQ6xgm1tbW
GZ5jxloidHCeJqqTP4s8F5c14r9nJZhid61ACyKgf3TmxgVVFZDXVr7Na/qfEcIb
GZeUXxQ3+VNKwjFf7MkSbjMTvEMOlnoqAX/cqP+CO/FoCW4xIOsbqsAikhehDQ0z
DUw0AHG69noZ/T9B1s7hZFaIIKr0NskRxNVPhCcrj8ILBq1zzdzbub/o1KsZg0FZ
kmK/hh7LIbp4Dj5fRKQQfoyQm1hHX40WJoGFUD4Mb27NMN8nf8bQKLcsn3B04A9B
CPbh+dLdbd+hzFclldy04O+WXznXt46cinJwPXZTzSUC9BMtSWJun0KwmVWYUuFO
8SIicNTmLw+sl0sUm2iPTZnBPtZK9IrsPetGGBr78mQ0gICT3bgz+mcXGw0dbSH2
xAs4rozrhvb5BHT0sLnDVQWNmFWqSpK/QbWnXpkzXtzmKRksqO00aM+USP5X9Y6w
VcHNgke7NCmX0VNXSAyFxeBHxuhoxCaoLUYVZPEvAKi9VPCdwiyNWTuXNQBm6Sx/
Jt6+zyu/CPsUE6QSjanQzULluC4vUapacPm2K1GDBPHwyZ1E5fqCjeswX2ZmuVr5
y7xgh4SjNBlLkugPzVoC046FlcknOHXxXPtRweTqG4bLgQHWLq/onJh6pZbfspNv
S6cUE2tb/8WAKvMenmDaYhdRJO0jXUah/U/qzxrT3yf26bPwM6zTESJL/mKUEVvi
RtIp0FvvS9LU4fCfk4ZShL+ItAFPg1VZ7sA2UK/J5sIGnmEfWNRbYL3sSh/Rrl1n
9Ny2rmX1VZMmGGdH0VMsGVtNvddCdZ+3M3kc1x/8tSTInW+ptEWkzBV87IimWLrk
TaO/noFuUnQhQG4ndWG3HYDZaofyKAjApmTNb4b/Lki671nbzb8OZiwMkhEBH83M
SQLEneBNjgekKISv4kX4G0ADHTbwNRIi4HXDKywsne2W0bl0Cte03au/XWb9U2Qo
EOZS5/wsFC/fRs+VR57o9sUNNQNoLvTxVj1X1oacla08fCqL4uwrNLLTLwR4JY5B
a03gO7noisbILhZNbkgZMevC60db6wd1IUDZ2jSbM0Ynb2FQbAvhgscCrA+7KckV
ts4RtvWwlC4vgJ5qywo45N4DO3nzXEbg1U457Zj8ugEg0uzpp5xAX9EmnRc3TYD2
ZYxI7H9RGOxia+xcYyQ3htXpRgZ8i4bGtrhcYEa65weHLO7s/Z0YJcBVJ2LC97sJ
EhG6NzRYmTyvOxDBTECfpGQrxYYy6Dgm9YnPo5aiAFuZ5/0MisXUa9td8NjLhMGn
0FtcPejm3SJMSFKPymvvlrYh4rqWwY7qr5q2qRzM5+U6q4+qvJ6YNe4h9nHcQd9M
HuRiO8dWpv4t1KyWmlubBttSEeiJj6AVxYz4bzTtL/60rwYf+Te9PX9etLT3EHLo
tANqzHiEvU9/Pn4MZA8guLc2ob4Eka5EBS6LIgmG713i0+egVYKEQ+xAAMAmr4H+
P/n2tJgxuZbBMhba/7ZVwCM79SaP6pxI3RnQ1abJInrk2atmcVP8j1aeE+8Gy9DX
JLLcatYhxo+rRBmtl+oByGoSs2axleAATZWVbU3Sq5JajpsEkehn1NDF6kqHSX97
eOX42v1Mi4JPFqkLtrBHjo1YxnNVML6XtHN42aYqFt5GcdjKRDQOlcHdGP7psPot
2LO2atE/jTKGg3j/BuAIu+/4APMauL9eqJaELfWop5oYHLxIFZmJHNcUoiZaHDJf
bja3s6lHwZ19M8bXtd8C7IPHXrRfs2l85tAbZOyZbZ53damrzpMaOTcwS+FpX9Dc
Th3hNLnpAB+75vH/LJkdTi4YNj1HIznpQJ87hVlpmAv/RHmqecFsUtqsCRDs6g5Y
FX0Zjhn/FHZotnab1GC4qLL3UDCC7aj5ZcbXKi/0Ewf+yw7wppxYgMZhxICI/BUo
4fIIjDLemPAgc5xnlQclpwvy4m9nJy7g6Xio1xxWXEOh0IkyHT23BdrhLlF1nqYy
8Nd6/8ubu2Sg8e5p29vVF8oLxANMvpymlw0QEiMy848dEdygPwRezMjuhLuaenxN
gyEmJlKzebymDlYfU5l6sqlMx9jqDU9DPgo+RjzLArgY4/Nbcu+Cb0JHQRp2zybo
3zn4K2/RLRMxPJlS83uxglPvKAOk3mov+6QRGvmH+t9J0myI0lQz3vgs9U7UcKzc
jwLn5fjm2oLdB5jH8/UHY86kXwBrvs7dYlSIDLgQNxkQWivYCulQdbsfbCvCsdI+
4o38kcRWUxrnA1WTmqTi8nR0tjrzan+4NGeeMJ3h7yLJq+updBXqfTfNp2ecKXGA
4yC5vMxcC/dLickGx1D4pLKIAbJKQ5YPEWG71lcloVxAPuDX6uuFdNyASnhtZ2m3
3V8Y2p0mTLfWS5J83LVVoCoemeWXp1Xy1UDMsLu5q48ZYZjUG61h5YQDrUvT556v
sWYwvDN6BC6umH3onG6ye5cbWo2X9Z0xPZ2mvSbw67LOWB592Sw4bFGwJx12ZdFd
E/wkBht0fEXnYeuIo5Td0sKIM3GHK7+JUTv+jRN/M+x+qHpWP8Mts4FTiTFV8NMj
+nTaqgt49Qz5Up6XsYmNOBFw91hNPAoCivnO9ZG9TBuD3bikqWPoBAzkdkBKXeUU
aEj2cNU4p83gPDXGlRsCYJe4Jk8RwguuM9ARGsgLfYU=
`protect END_PROTECTED
