`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bjdKWv8kbo5fak8110nqzqeHwm2lTLhjI+HLD5YvsK3Q2+aBFtDeheF2Aejneax7
DFxg0JVDXRJIfaGvTNx2L5pWStNyqT74TIilcHzVTsfIqPksl4FZsIc6Ub8wl+u0
h5DGG/v8oAtwjp6GcU6aXb5BUS1uxMyCkceIMmAx4WqmWYwe/pZE2dk/qvRI9aDJ
EwswzcFAgb6opDAAgWxZrlD8UzHhB011sm1nc9YstPyzJs9Esg4F+MEGNhHQIv4n
5Pt0N0kaz1BodfT2/HNaGzTJkV5J06CA/3HqnkdmP7ODZ8fUJXL0BRqTMbvZz8Wt
HHGKOuWsIof0458aJzGQUvNf6ir4KV0wJKiJeDf3SIc=
`protect END_PROTECTED
