`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
KHqbzjNDfyunY/s59BtMEoL1NcabrOHUziKmSp9507wpk1TM58j0b+xUukksow6k
u4YQnbycpdux1YeZSbYz3KK+r5RPPA6cDct4USBW5+LPevK3bRL6Jh/rbosdmRyO
fA3afL/+0eRn3mY7kr7aKH7QsbrIWGPig/urBF8nRHqwXPTSBNymkHuf/A8Aq8K8
qs0WEj6u+sVWC+mfjdpXS9yfcKDTaWKSarjBT0ab8BiDolXsnqYI/zIEDHMDwK2N
31tQOTGNqwYnCVtZ0zexy3p2cQtfQ4Bi8OFGoeSqspoEoHInPoZTg2TdBKyPpfl8
abS35kjHIku8eahelewCeBf9SJhXXAL4torbSxwH5fRM2G4XY9f87nUYEQ2Xihwa
MKz+EPYxUvc1W/qXNMRU3sKDbiaAkzXyYsXc5BQOnfo=
`protect END_PROTECTED
