`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGDwWRtgykwWCJ3LRUTdzuPzh2ARfHJIvHYLxCgQTTgR
9acKWT6ETE2+030jfosO/Jfj2ndAtOvpGrwBOGDBteeBXAiASJtHVusw6EGkDJqv
CyuSUvJbks8LhgWfogl9sO30NvJGJv01vJvEfOtV7HUO43BBMBCgTwUsCKPiK5Of
u/Y0OU7WzgysBYyiXMoilh5tZc6RGVfShoRXlvnXBiKgHup1oOmn6REneX1LqJtT
0Q5UsV6EZL/OWV9vKHl0IB0GX5dYVoFOCWjCFOwcwhdEPR+Q/2rEpq49Y0ROy7ZC
q4lZ59NacJxu/QC6hUBMk4iXp5YXRAQIa3StIUZv8VOX0DgF6m/IvFQvKi5qG5dd
95+qnOKLeX+Q/kZD4bAiFZnWecsvG6T59hEPKkKEMK82J78GtfdNQ9SI50Oen+o2
Sz2uWYmPwRQCXhfk6wDoPlNyRq3arhyDBeyDtlpK9MK9TjLmPd46qD2kAgtOCODw
PX5Do8FV5+t0TdYtPB7RZc4kMnAqxm3jYA0Q6esenDwqCaXXLjIVNZPC/lk5xBV9
`protect END_PROTECTED
