`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abT2z4vAu1InoixeAjOi6m7raGBSsgAf2R0aeFXZwFEt
p6guHtX9MwMGgzTZKgTyt2FVoAe6mIphXZdZMYmJfhQW567RYv/4oxADfdnY2kkO
HLa1CPbDcgsD9qDpbQRXKH3VPEwbcOtDBqZlpxoZsNETpk5lBlKfdEntws2rEm7y
YVoYR1L1867ZhbYGfG9+Ufn+lrjtu1dfDbox0CTcMnDLWTmLMSZxLH03/4zmNqeM
MxoYGUoCaOTp0VezRV54Kux14etPQRCvJa5yPvrfdwXuMzfkzur+/8Cudi9tdhbr
UJIqzLBC+u5QNBkIhc6rnzGwNBRyr2l1uy4oMerLvP7EpIAqn4qUf5HpLDnsC8A0
IcOpf2F+tyUryNfDBGYWMEqkEZC7/rhQUHVaqYU8+ZFeuFxgoc0IjWVg3S2KoWQx
WTXYxpWaKZ+22RtfiL0zZQZNdbCbIqnZ7ieyTAPWKE7chCl0BhUBwPZjpmCkDLAd
W8uo53RemrHWQlaQu94327g/myWf/tQ3Ix3/LYt+Mp17dl/CoPDJXaEPtMxTX3Bv
QqbfErVNw/Uh6zdLZXFMPcgfysXnmB7xXzs0gAf9ldSItqdYTsLSoBRAkPhvkBkF
JEB+ipZJzFUsWCgrVYCsedPQ5lZsnoqRiZOkS6tv1MSIjJYPl+eSi9VGAAkMLtba
7EG5BscP802/6meoSiLddRq4SfpiPGd3KAjqKr977COHm0jIcc2NrjQpxDchXmbu
/k0r/nnHrA9I2VSLW3s0dScFN8z4MfSjEKBrNIqdVr3pX4IbcirOcbyVMoNcsRLS
RT+gRX98+AnG5lt9UlGFjlqbhj0mVeFnj+H4Rcla/mLOZLlL/4v9CLKm7Bw4Y0Dc
247zKZUzdO40QZarC+n2yk0qImWBXvCslmoyGlf7sXfpKiSOi4fHfU+rLANa79LF
CTkhHJBCGaFCYQc3HYRMOkcG6rwEJHOLMVZ6ugRoS/kciVxJqatyzHNfPmWH4cGm
MRq9/ydIO5J4lpaJCbnOCrHu97d6STUIv0AzM4lCj3V3CrL4BTcKu+apHAaG9QR1
BqotHeQ5CqhgyJ8Fj6TC98+M46u4QJ9Juk09qb9VHUJu1EZNSF6pL863mdtriKir
HozagVbABD2ngMMj3wnla4goB5ayWw7Q2jRc8c22Ihz6+YT5JMXI3Yb8M9sShh5T
0IN72pgHCceW9wyNbR/nsviMlkIA4cfY13Lf7nIB2+5lrn6rFCDGNSx+R3ZacENY
Xjc5HTjKmGAwaHtT1+r3Hwd1jH7fi9eAJh2rmv7+2+w8y5vlJ4Yq69cI3QzBZxuj
02bSkVkJyboOFhKpHsNwbaC6jP15aQuvoOBXuXO0YMRUB/nmjXeYXhqSs7CRvY3W
tDC7nxkaK0V+ldBz6UffbuuTy7Q9uIvFRGz2I/K5DmKN4I9h2gO62KzlcrdBtyL2
vFxDhrCkyYCJYqezYVY4L1bvAZSaT01nYEaot0NfnAvZYePxxaneQZ2ZyqftJL+f
pvLpH8vJ3i4DhlQpLZZmUqahitFJlBxUcxzpnIdMrCfM3nA+qOdEJp4ZRBg3ZbTE
+EKFD4jimV8G5cyMZ0i9mu0DSeWRsbL/5n5kDEvNXOSMnIreoiQccxatp/KF5cOr
DEURIQZRVvLEUpdC8upACjkwBeMsuwbU2nffVO+MGiXCOE1vMr3LfP16/sr58vCF
cq4IdSh01GhbKHjhZEzq8A9iphCpfYZqNFSxTVdQrh9h8xoOpz48pOq3xL+ErghH
u6G9k4W86kWEla5CGd5sh+FCJzT4NnM3xgchPBc6KKdwMo2z0h5EWsJqVmR1mt3o
8sohCF/U/VvlAJme5IzgLleYhGYvhQfyEQ+nj0+xRh7sGVBQ7yTTHublgg4F+EL6
Do1QHn+mDQSvD07zi4/aZNP15hKILkE+w5RmJ5VFbGS+VuR/ySFS/ZKBf5npzIYJ
rZ6OjsRKXVwIdi4vgAN94RRpXcegU6zfzkb1nK68rFNyPhgsw/IwsvoUI7LNzhDW
PiHVEYu1EKVFp5x4nQiAZnSl9G9TNiSjf29WMxdAiDCG/d1Us9rjAJtXzR8M4eTN
SZxPhTbhbEgWckbd0D3rtAte4P3MTQPD4gU5TXOJ+V52J/R6TCUOQNzvKlwDacdn
TqiuASVAxfm8f8DFwVCFMCJjF8/4sRGMXExeRUF/OL9KZP0MOsNUrRN7rXJ/QTEz
bLV7uua1TjwzrGWM2d8/tfHhSXgoPAvFiet9mfV37FJNikI7zGcghzRELWrMwYST
JlHDBiEZt9LTxrCPNdsZIT/YXSPHx2P98AkpkTrvBrdbW78CO6nud7gZLOfatygb
JLuB6JjVJQLKwQSNjzuX86QuZUcNzJYtTQF6d02LMMGs5siiwON8Eue/n1WkoLPh
Mw6PcP3nImMVuc/ySgi9gp1yc3D3W7sJ78qZLV+Jg7x506GhplFYeYpROsNYN0tl
lAlCzadziqrcdHXjgux5Y/e2nBStxSW6OPwUOQEDAGbSPWcXcTxkHY4mDXN0uxbk
4dnLy4vBfkXixLSrLwUIzezlqCjlJ4kyR0pP1uWq9AUKzM/IxluPJDMOWsbPnRC9
Yr04kN0DQURG1G+Pthd0bNGEnkfV3B5xsIFB577MtpcwRDOcgZSS/c9pQWJlMhgm
hEkFURRuKj3ja+iWAmETYTZciz3mrlGbv4C6nwSfiOsijrr4y4blsh0mrKmnytUa
sgWPdH+wdaV9UwYwIe+CFCLTs94xp/v9TQhAoA/pDFMwtgRH5Dc5BC2s559LSCaL
XED4LO/BwJRm/QeGnEsa5l91VJC0/uEi4OBdzdcMfoYNw6TuCMIlb6jdFRcEv63D
b/xbV/hZK64Co0JygrYHsrXvcFxk6MikHGWjDz0I/M3bFLjd33opeZpqgRsSfpaO
XxWFLDqzxegguOCq2R0m10MUDsEEQ/zrpoRZNVY+hQZn37ab2bBPKvZIQdIjLw9e
rwHcNN8n/gmBsjbbSZjX1NpLpTkCDw4XBzWJuRIqFAXW8njW9jhKra1YISblvccv
C6H2o9wvkavYi6FwxuXgScxLHhhhd3pdoUUzSTmRhnTCjLMuR6aU48GmzxJgWXm+
Ax1YohXS9tZ6FxXZJKwOT+GYG0X0XHjAb51c6v83v/G473o4uFmyTitaZ7uxigE+
fjpN15/V3SmYFALJIPsavoFuE78SgPkTEQe8YWr4t5r+GVH8SwepuOBzhKGOBHaj
dzgrclXFAxHHx8qabxr1S6rbe8Oo6WTzJVK+TLMuT7KaigUMAZoat1cVvaGc9B91
s3cmRCvntJo1wjHkuaa2b78vWf+pc8AA6vzg+AiMmMuWfB8CpR+VHXXtnNQhWY5E
M560TGn8ylys/qJUND0+K6mjgsTqDr9O3Tnh4iYZy1GT4zCpN+ozcxcKDJjfSvn6
t3ubXuHSBCJIBHrO+0U3Eai+YScDpmUYiO1X2Uss3KopyR++rtt++HkkZfyB+fGW
8pq/h8YPR27pRZMtFGV0Wa3QTP+15ZzhGmHfQbzT7yEJKerzQNqJJA0nP5MFE0rv
5gGd7kYcFRB8d8gazWvW2Fl0M8oSY47A2YE06TXeAWx5Q2/ple+l39Bo/uEpz7+e
MpYrcKs/8IVnbsThXQ8U+YHMimQqBMkujHrXMNTA5U7a9jVpKkoNWGJEIFEMFkKo
LPUBfdthedI4EF09PCixtMkoxmtn4GC+tFF07txpSNvSYRHpFPHBpraBqZ3t2btZ
kk8AaRW8738sbc1F/O9O93/6wbliP+Ykks40j2wD2UiPP8d7BlrjaWqNNtKvntE6
oleOxi/UUFTC+veMh/29u3XLjw/9XcKwG920aaUfWwW3gkGKSBQtcD/skN7fFAoT
k9blE/eASfXyG/I97EEPjXHvaYUeTWVZsQrTblSo61onMNfKLD0yfYf/vMsSsuik
tollPW5Mz5fp7ZP+c6dKgyUt97oLxfHlOXnydznhFiIIoUheFiOsE8BbPIUllPSC
iVpOT3KXOXnRi6bzzImu0pFO0k87Q3uKgHNBd/Jkr9h+WEoQAbhkPUsSzSO2iWGy
sN4ErpowLiRkzhPyOmqSFGLVcUSuUCuHfxQ98210LAUzHXKVwCnwbAcfRe72NWsb
NTtJnAGEwbV/pva4MQErOdXuTVlnH6prC8N2JdVOA0P+BPgebLde5lzWEoRrXpzf
+YA54N1zDhPE2nhCzoKAgVtR3Fj3hYf8dr7+ufKcJY/tSGWB1zth1w6wyOGpJtna
s44j660JDjYUj1AP39QqbjAqKk214b+OnTyxgm0/h54JLhEwZ5VT2KuAW92tagen
+VxXk4iYj7YotZUi1GCEcFM7DsP1IUTNtsZdfmEXGUzqG0bchKHw6Czc5pOwtqCH
NUY2sghgf9sxUUZ+qls8gxHBcv2kIeNaxcqcSmnENgyDtKDJEYHxzmgQVPGrSfVK
jeRVE2vzRFE9exNeoWEitvCvRrTkMScVsmQggSZalj3YLhD+UYEiY8mmS21vS987
48BEKHNTdA8ks+OsshAmrdFEVw/PCirbgDsWpiIJ+bvPVSfwmH8lvhpAqWCzBVBS
QqvsO2U4O59SMV0YIIJZDd3G0qGQ1TiDeA6Z6keK/Ro0glcg+anNjtWJ/r0QEdJo
sQLtowmm7y5C1w67hsbCMCbRSlV1cDF+U0JAfqf8IHsIuOTbOLmQOyLEyx4cnymZ
kTsXLAX168szCSgAmXdpVg+c38RpSkE/ItVvHDTaHiKUbqqAh3NeZfxxq5PaZYDR
hMtURjTzkU8LdqVJ0r/gzlFVX4BHsvEknU0q0gFNYjD6ankwI6GkDoBqameO9pSg
9rB8llAbmtKzEZc7LQrY/L/lusZrF5AGWZJnZDAoJMZIJp3LTrSQMF5pKCOGc84V
x/SinLfLof0j/J3JZqc0+vOgktm4J1TsS3WyFGeLm2MJjH3hprS8Ijqh5mHkVVjm
uNQ/ZqxI7YBTNP+8hs35BVn9A99RNeal5zZS7s7dOC+BMNdCCPnwx+apSX6uGM6n
+yG89J64PA+JhEPMkzD/nZg+IZNqz0Ud57njUvL+YA5u4J1UyNujXNLlSqFIHwq3
JoYySIRSE1Fzdc6B/GDyD3SuuFVtnhWGPrkrByT8oub/gfV9khjie/f24b1vz2Rd
bsINngvXa2HnV8+Y+jl6y3TRad4dGtbPt1dB1NuHcMhQ38W2wBOLB2UguxrYdkZ2
XKGu/OtAYgdlm9A1lwHzpHCpvsChj6jeEl/sMWgd75gxoTS1ZHNJumYl/P1Yhdlb
KPkEPSNa0pjbDMGR3Qy/YVRA+DUzQanUeiF1OgH+MQm9gNWf8/GZACF8hDxBrw5B
va4SBGXpgGC5J+NYCJnIyODAEb+ZsgP6KqYmCM782upUT70WQjxX805CiMb2EwQa
hrGfjk36ITX2+5T1Qxd4o6cLd3qY6JsO1IgLx8pWghQeJGQue4ztf5DIvsqpEGe/
Zkq2MB8O5n32fymH1OZno7HGnB7G6d5kkJ81edcZ7aWFhGvzNm+etglra14dHisF
8Y3vmNzrLQyuXzGKEe21Xnsh5yKc3iwsLcCH3O5zGxfAsu934b2yBnIXINm36++t
bG+aZxFFa7rv8UN00bIgZMSE5VKgfMp17jkgLwdwcFXvJkRvLKE8g7BOgVKGajNs
Bxh8fi5Fk1NC1zaacHoPFKHa1bN1koB/+XkIOZs9eHWlwhQ6xcPGiHATT/3WGEAC
06kNe2q/bqwaGy310c71ohv2QRFbZfIKmr34fIBy3YyGF6uV4qP25jE2vhvQKme7
EwTjMHrU0Kf7lzmXTVdCKDXsACmo8ubcMli3UheTkVzTu/ys8yCqw1HFmAe4iU4h
zHZiBFKGBKt6RGKMecYfkgutP0fk4yhn6d2AE8ITVa4TBvyYlE9MGp95Be0eA8cM
MfX/RpCuFijzbpQObttKYjzJoFho2KqaEPyIMW1+JQmJzuaw1inQcb4XRqE7mYzW
Qh2LzKAqS2C6v0C0b729A4b79//BBa8CEW2yg14aQtR2YvPQr7zVAzSpz6bvOop3
hEHxG1plJ6YzRJrJyXgfoZRYU72NK3FRGQ11G1UpuKsCjGa86+sm4FW6mPuMnvVX
ng9Sy7Exu6dmtxKK0j6C97lZwVIWqBZjxGIquvj/pfo4s3p3Xr+9Hn1KuPOelNb+
ldmmSUXspMDlx1PDbwk4xVqW99m7JpscrjJEhtSspOP/uY4JYBrOCj8wdlEqPVfs
Uiom8ftgPo9/IElptMIm/ECLdLFq23HUYEE4fJSqhPmxd6KFfCBk8JSTMLkMvfkE
fK5t9bzuWaaLsJDnMDTKdyi9IOJL9KgM4JMOxrat9Yqs9gbB11KXeLiK391uH4We
WHK2q//c6GNP8M1hK19dHF9DaMMB+1+gjKkjVxAU1jii9kruPcGOHF/dzXTAjDCi
SwoHfs3wQnme+veeiiqdHkA2V31rSBdEmcuKgf23umfm1wiqoDPLWWsK+izx2j6R
Zwx2Wxs6Hn6l51Z9IUDuLH01E6qJJ+vqKZf9ifa4uBNrLOTZcMq12hfg6AtmbabC
drHDXCcjd5Q2ZJzD5u8sr/C/N87v8J/epESWurDfBMa4TLbN9RPBZmHXNY3GKEFQ
RX7awAAhj6UA8Ahh03kdUKpRedsFTIiM+NF+l9XHJcbC1ysOMFdUQ3Rvo3ZQasCN
zDN+aV9hHvNnRXlOhLWCjW4WmLpk/LjpXuLWtDv3LxJPOVeQxiXTphpOuYRyzBon
pGdSyL03hN5LubucJqIRVer/CfkOr7bKDP57PpYtMXVI8e0F1xXEO1Jf4ui+IfS1
Ebbe2qnEeuZuGKdccdnVRqqxZQcC/4jOpiBS2Nl1DnsJsPlk9cxLH7TpPD8acCLO
n7+P7oi6szf2ZetIJSEUWx/OSXqxzj+i6lnruhn7qJVD5c6HonBKBU7HV96/aDcY
CDXpE5mFTqkpXxLkgXzqjK5NVzY07LrOPd8DZ/cmv1zoDxqWhHLHLgT9B7vTBCXW
YSaKRn4w4u7+cUQng9o8Ic8QmlqSHnUjVf6cPTDeHSvVOSpM8tu4yTor4vmu52DL
gfBSSgeexyoBd55f9k8P7iFjr+A4YKi0o+5Lnj149BZa5IllLUHNHvcli97gPyXJ
ZTndc33B1alnv2qi9FwWHrEVtCp1xLqb01/vP6wO7rIH0F5yGI8/bYUtUTZ1flcD
GOSsup6FEccKTWyHMPcNXtu/zT4wbNX/cd5qxOhUHTj0MEDtWqtwSLM0qv2a4SPO
3k+j8TT/Faolz0IBKKUZ2nN1QEbLz4OCBKN/ciZZ5MOgmdKoAQ5LhCns+/mSQzru
KENZ9NRUAnL3yQAI0K96NHt0VfSgWwcNeSB3em0SFBM8uc1qcMTFtzCrlHb3ua5m
eG/OVRatmMNpXK5L0CwOogHUExgii91nJg51WN4/lzgkxhQoUbHSUqLEZMIzyaIu
GAUfOv8XRoxc14/NFwSzkO9c9K2jGXVgxzbthBWWcux5fP1WnDr9qgvX8x79YLGM
JeNYb1eWjXaWycQNAM2u0GCQ1bn8FB6DAZTpxXSC2/HDZ7fqu0UDa2+hKn7rvGdc
G65t0wSM422jgBnu4AhddY/TZMwIKO5+7SSln7LJnOi4oLBuH+wi9+w4yewiOPvD
oBSb0KcCL6+j+8Iv+huejCmKF6WeaG5DTrtXLJKrq1dhMZ9CZ0nK/N28+l6bU8l6
mWURsKQwz8RB/dsgPbs7YTTPe/mmQ5nnVzs5yLzwlQicc2YokhlLTEmoABWzGEne
vjW6lpjiJtQRcsmN2srfnTSxgVdrURhOhwwM6QgsDIK6094yBU2I3TCC32UI95KO
amImUOzVUmtAYtVly2KnGEETxEF4YZZgDDzd0mK63VSq26Sqwku9AW1SEheIx+kN
dSz/tvWAg0bhFT5l/I8wNdGgHAA3DCYm6ePsR3qyw53aoQYCHYIwzFm/z6NxMJVo
3nYO+UrOszRH6CjT62IBCTDryRofTclB3avdVn84jW8AKkFfagEpAgoYGblwrkkv
tE1A0h3YU7R18fBI/GiY2iKxoxi2d3SWI8CTv6jU+ADBYl5oA2PVOStqu51ZllN6
OaQfgCGkW83hc3KYt1vilNDjOOct9wK5uUHM6U+FDmUDSAQ18BMnorQC3YW+7oj3
3sbyBgQBlCh32Gjipyv2/Ng3aGTQ2tUTAAuI+vfCBsMHfAqkQAl7WcxFQ4T4r1hf
zjjbrZ740V1CI39Q5xqjwCS1d2fXbyJVRutpyN7Hx7nmcM1rNrbMIWLG0YsjqzBs
7BxOqMPP09Xf8ouCQqoRx1qcNuwJEOJhbIwGWhTmhlSnirOtoInIaulC8WYBOMvG
zx6XIQr7oK4L+CnWekZhH/NdtI8rHa4TCxYC9nrsI/N1xlsOLxJFNI1PGCXEuY/Z
8nsGU1FCq6qzEyvhGrsL1cETE7g/YGvj87RrrfZYf3PsuxrpTijKJaGBPgMzDVt0
flNiruauFJC2IUe5VKeBWTjG2qHj0zFuCbh5y1xmi52WWASGXrJSXX5Nyh4UyY6s
JEstuf7pv5bAwKN/cuUCKSeDSeFAU9WdN1SLAFh71xNVUtUhTUbSzQ1uCDv5cidf
J+VwVZA+9OmUc6UWeBGuJlKh7NAMRMxMdcBhGSWxZFOvfACDXcrtORkJIIxJ7nNt
xZeJXdA7zo+Eoyf8hkoSSZuEt2HMTfYlPJcAMxPs+gjUAXykDwL6PPlaKXN1ljKh
VG65nPaT2S9YSmE0C21u/sMOxYQQFfIzHrpXt5QmdYylG4bjph5vX680KCt+Ll3s
H7lzsahPpR30RRuvhnJ0gmo2b1/ze3FME/FSp37UB3OrOPySYyMeXM7KHEjDUKS+
L9t/njQPWQGSblyyWp1pWTJAIVQVzSiDvBAgFJTZ42BBcDctq/d6IAS4stZjV56t
nIpsFgluulTToR0d8SrMvwAlWMF3eKFOLCg+kUpDS1zY3MUcGGNT2E646glDitt5
+UXk5GMSOYwHsuwdNgsASF+6YYQKZsgkybLmRKepnqcRPWxo5/aFwJQZKXpg34hd
GZkzzzPmuEUyHAh+F8lkxPQKinrjHzsu6F7EZSgzsCC0IqKPsbUjj5cywZsSZ0+5
qTYmqIJagix+0Hy25gGjuQcgtLRpY7xpInNuTdtCKHDBhXXg3jPh8/iCa9m8QiLJ
JbaxoIEtfPo+0+JE7qYc2R8bOWslcISSURH4BcFRfllFJmNxXsXD0wvahJ4x9KGm
GnGeoDgHrzn/zH7rWIj9Lvg/bU60zVTq8DqA4xqllIwhIYbZ0/q/zQc5oI04r8R1
qH5ioxvQMRmH0m703AKb3NgzomC4mhUumkgCYPk9Ao+lM38cKbiIJWGGnu8WU9h8
IAF4M8/BzpevmcsYj74yKmd+OEmNnGkZm2cXk0z1s0ciNbcSqbYQ5hdMG40ir7E+
mgcqkj44K+FYs/CC8UimkY64tw91g5x0aYj3thqOpdwRhozVVhWmDzxh7eJfhD1d
0BYwIrOaEi71NqbcwnDcLz4D8/4ppKfonaFdd5ooSYhH0j3OYaforxunOmGXpvYD
fhuTILQSuJdH3yZ/r+b7f68h26S2V3UpLrJcrRrihdY7MCHrOujHchH8fjoIfBv/
GnMBtcbStglwtWQmWdhdxZJH8qykFNNP2xpiOIng6dlAKhqCiejl7ujTa1n3dquj
FaJbnDU9jFiXCYjDUlZqMgInYEs3NwYDpvpMtfR6+SplBfwl3hDMol7/m/etqKtN
e0GVIRabWNQW46C72y0ZCYb6ZZItwgAVA2haIiBn2wQw4LXin1zajPHCawsvOkm6
DyTdJKasIbVzoIbShG8n07XIRhRRomcwK3zKLtENFbQa4OjUQ9FM53kihg4Chlsf
piTPPxVLjBSCn8K611MZC07DuXHWD+ZXKar9f0cF6rEmAlC0W9wQUHA/QqmFOFSH
Z1psvaMrGN8+OrMerzUpplLWwzW7IZdYMpgljBWsQPHLCQmzwpwfiSkf8sBwqffb
k6pRnrTZ/HStyCugIthvyJ4VWsRRA+8CbAuTdFkl3klQNNgrs0f9xM+fnOy0AJAr
lcMNA+mIdoI9j37HZUC4oYrFJWCjaYYO6uHzrnzB9xszUxUt5kuJ3nG+RhXqnO6q
iYCEiPYmByNTvh+FGI46ZMtV1/89lc5UHaLqOfe1LxQ5a9m3ZXPKlKVhNWROiSIe
ex6AP8GwOQ3UA+v0pqKZLRMhlaNafh52b8Z2TXUAeZJ+kflP3tm3RsTI+CDehz21
VZB/9xTQaspm3GiUsbHvRa6BEfe95ZS09BDvQQGvR2G9UZ1O0llUtraEX5bUzZ+S
TJe4mROYcvKxw3E4PKgOc8A+RwE05FgCH8KKc0iCrEpltN32h54O6Bg0aCnQzCW2
RVIus8fU+C/K78bxPEO5ELHllkSd4JfY2gC6XlGS6KF+FOUQW6Rroluwx+3UYsYH
leU5NBXzsvRbtkkR6md6aUyRupLK0Pc4waxHj66wuT0WtahltwZVBbSOfupWmOpG
5mykK2XlbLTeWjB/SB7yYALyvuyeorQjyAfRtmYnMkHlCS196gOTgtsAkxTIbgHm
Bl6CxwXchQA6YB+OcNhYDz0HXMAYumhq9k/QT/z0ectE9tF86cnfe08wFOeFjGUd
xeo+kFilaO1S8LSHWRXGLe2MJ263LVrMDUyojvbQsnOQCXIqRn4phw25megKkfBH
+e6utoBSt/LMGKgxW8KM0x8iZTGdA13Lazj12Y6aitj4yODb7/qrcMADXzl/9o3Z
yIUagnZHSnrZKzBTDT61t23nqaQs+gVMRX5/RGI+6dtD633MrmH8Upssp23kBNVS
lTGar9OAT3V8xgqgx3n4yMQsgt5zjIRaghl6I8xyd8/kyhb571ZKNhbaMByaVZuP
k3m+sVOOscuoPjXwo1z5u2UXXPYnJCxR9bCgtFgIXdayboH/rMnsgJ+Ho6iuvB76
ml1HFvME69ATzfPoyaM6WgsK8r87KHoCyKXXwnS083GN8eZDWrr0wm0/gI2ITZNi
bL8VGIInZHWVhzIXRcWWr++tM3Ui7gy7Lx7jL87s+R1f+P3hYFhRT9Hqs7DjL96g
wd77yuypd+Wh34CZb+Gd1q9ja3LhqSVnqmihVM1gNwiVSgLnm0B4DSOMETP2BcWK
u3K7op9dahZVJK+lJ+wPj2R5T4fcsgKbLNcF9zM8osJqppQHO/U4VfF3Apo4TbDy
vurnyaFpbqm7RDcyfGL+MMmZOWRSOeCuKgH8ynOW3SIjCjpPF6UGCValWeAmTWhA
HjO+7/TSwBm7E5AEGk/ooJnm5jyVOQT6eYR1SvGmjmKc9YPykVxL5fosgjYIIILK
HReEIOyeqoA9/WTtCd6f5CXWX61OZbnUnG5xc4IbVZSd7csyAocfuMXsTSGbOkjz
8OTqdmnnCaH9/KpxgRif5LrMLLY8HXjvsUOVdORdjoKRStjuslLL9wdL4i+xt38b
UpTjFpTuME4Do5ykLjscBIoZblt/VX5EKeHVWfZ2GU9B5L6OvASEa0Izeq1OmxF4
QlnjMFFZ8S7FafzxJRF3fmq9ZarCx90kQs6P4Bi6fY/NT8gAje3ViT87Jwan4uNc
K0Hs0YDcAJcI6CetvBUcZVyn53X2MOmtyBmvzJSzcBWkQhtGRoYTeA+2M3RLlcXW
VIRUG5+iI0gLWfBjzr6k9E8tzcFu4ReRPwcv4BE5nYi02ORFwS1IbwBeFx6lAwT0
VMaN3VTz1D64N4qsBxu23YW8JgzLu77ovLLw+H71zatOSG0Dlhb2lrei42Bgpmdw
RyecR4kN0MiealcbNqvh2Qre2T4qHQ1z3Lh172vF1jth1DosN4Lx14WuwRiMEKVo
J3j8E1WzpzpBHKotC6SJBANOw2cP3Ijfc80qCied3QADr5HUFFYUmuPvRkEkclFa
o1uiAkNeWlEN+KlvX2ko6o/VgZ1Yq2F2PEkLiRyCxpIpfrnGEnNBO3LzmY/Jar05
XXpFUNfPofJ0BHU+F4AkmPjqOKGtDrljHcXoXl6uHmkRO7gZsPVD1wBfMKw5Gcvt
7t9ROdunsiJXcZq5P3rbFFMXxaytqPUSeiHl8L3EKZ9uHMoiUCld99SxQRKbLO1X
jHyeFVn5MPJ1ZjKhq+OVhqCD5ak6LTWf9BbThVUJEMTTfE4Vyjtn/HyThCgN77ry
Dbc8tXGItdpLbrzSbIkqCjey0181KeX9CPCCvedAB0hYn4Xq3kV1mEagCTE5og8O
3ihv3ja3bEj3BneDK0+Mr5IunCVjyt2DmZdqk3hO/zDxm/aTp+1x/CNZk/4QdYLM
dhzvTrTtBMlzdmJlfHm3ddoWEdOTgBzBM6PvQYUhWYHLvp/F4ykBv0l/JMLwbCNk
hCCqLfVNzqrDe1FyZSs5LyzuUGFxZo40PPU3OP0qUua/AAvPg8wOoxkvtH227vE8
NrAin3GV0KVzErDzV+liCflGp9V/W4N3OPyQmNb5tfdgWvgijWkvB0V7+62KDkwR
oo/ROKkb6g4pc0BFXwjZstymoZsG5CptGnStPaSm/KZPPqpp1CaA6UapswegP7TT
7hbBO8E+5d26rY0AOmdIrhERDRI8ZMpXmiAWW4gWUzOOFH0rp62azdho1vn44Cm0
ikZoEe6MYQO5BmG7Hd3Q2o8P3JTn2TdGcfJkNDj5k585dvIgNsrCMvxtWpaoiGMN
lvWf6aln3PGLP1WHAV5Kc3/Bh0GRFZ1wncSktK7Z+/mYPlJpXKzxBCF3xHlccUJ7
KT0eOXGjdVlg2FkdlslMDb2UlKaAAy1gUyZlyWTLpuLZWbwG3FfXdpzGvD5Ymzkn
3Yfsco4J9+fF3X+egW9XnVbttVzBnWluMis/ZOzxZkbxV1ucCXufVkE98lVKemvg
Nz+sYqEsq3WVtHtbsNVj1Uf6g1cIo1BW1XWom2nhJKqwTU+ZMTAV584FW4eKnuUY
NGiaT90XNlxJnL7j7O+pQVp6+dbrAzgMCSifYJy+wiynEkNXhSKHN2SMgUppm6dy
IgESqgB1gpLWAl8W+rO6LQi0ldDlXMAIKFnMPo15ybuvSCAvL5WU9VyfLd8/PP4q
RiEbl3OlRgtoJCivNI0Ir+zessIgX7vC+qctBZDcD7hdXpDHOEDUM15pKZUcfzTR
M2jvUlPiY+S0JS+0XS4UrqAs4DUoTey4RJbIUg11bEZHSyhPMYO8cM+TFlRoJ3kd
R0xNoXcSvHb3yjSOTrVxamcABER00gs9yWHZIXLrBEOsZ+Us78tvcnIbS0vuuq4p
dc1uAdNCbRHLn5OnBquzVEQgJuKQQeUNZb1o4GV/ahFQKf/uPuXgszJE2zlU0u86
tYLNStcoIa4/UHRGVf5x6g/mOeDR/x2hRivbwF34CLlBuRq9ur8C7CR4hHCVJ2cO
DmRPv9WLCeq6fn6i2zdcoigB3d6iP8jqIdwGMzP/KNsynJDiEFZhtTgaVKhtUoLq
PKJBB7Gp2FxscdTAR/A253X0HjPiU0IqWpUm94QDpCu3vvtKM2QpI1qs2H22srPf
NOKS9wUfgomfB5n7cLkNYG5jFtNT/xZNCXCDt3QcRCklnco8yrgOHBfDqihSC+v3
hhWYyuVnR392LfO/+xPCpRDqNi+gWLJTaHy/eafi8/c5nbZx8jWNd2K3KJtkyXqq
7/9fwnvcyMxe3WLH/x1JaHPu2k3iVwzhrOo7ghAGqefoUV8q3GphTSDJCC0gR0oL
674rY98MwE1BboHoMYfYMW4/MSw0AMITUhYP3zX1woE6FBETShDOM6vRzudchxgB
5Rwd/17X8230zpEz5FcvxBYR2q1fRdPexYcyLb8sN9UaxiMFnTQPA2CwqhCuZnTd
OYUMPFUUZSRuWOPfxUo8D2J+fin1wHGNhZ8JT2Rj4ztWBpD9m86RvuSE+o2SGIzf
OJxpC6jm23ieqWZ1/Oaba8HXFtboyxKpJjM+dzvv9v2BsAxPIzUPeadSech4CD8Z
ijOG6Z7OpJb1qgy0qL0HxLwlLNshWTZ5Ji0qShppWV9udIhgadhpm4u4BNgEtZHM
PzgBZKfu5iZSNh3CFqR2MQpCDa9sIAP6HBTUB6uq8Sl0JyGIVEUPlREX3/hP+fmd
IhWDelp7aKn2hJP0SeAwuCFBaLZkJp+8UxU96tTRHytlH2/ld8HuOWTfxNznhvIa
KHX14y0y4Fio+d9v7WufWrf5xibm5yu4hUstWivCU/qdutBxtcvhpZjP+PMzMRiY
s+Cp/lr+5y9Pp/pXkXmdsLnaZQ3ebabZcmi0ccZeTtAw6qMdoQIwEJE72Y9tpqRu
VJiPgw1GpAHr8ybdap2BQJ0KiyH5spKaI3w/Cc+lF0aIsZB3PsT9VafjNhPY2Nkr
oWj79I4i2b/UqiWr5DtLNo+78Wwgf2688OIp/l0OpqzhmGxsYjlrYc7dVj29zETW
zXd6tSV5hhor+4OHdm+Tc0Z24NNRvjN10RkT5b7U53Sl1f0Kj8veTEgmONeGnt6G
5oyyw0nDDXWZU6PRAldJM2Xae4WKmK87snZqH+pOKGC4BKLw83VqZeKmpkRrVuPp
/2uvJ24Ddv1ZnkU2TuRrMJWPyfF2BpqYwspUdlRvxzgtiyY4GqBqaV2HZzseXgvP
P+2viLzXFrtLTswOwBm0mej9tcIN0qDqvTT15uYAE0/WH6AbPKN32Xp2Yh+CwTA/
lqwYmYoXnSLuFt2PRkafphTD+f5pJJGC9raYOCNYgWu/N21b2Ng/NMMQSgTlUqXG
tSegoeCDWseOHYmGdEnqlivB82/iQc508erZw+sg373/C5x1OgNoJrUfD39Kfixw
tb4HSbhh1EfjvQKb9NVceKKUv0bHf+H3rgc6dFCZv6h4lImGu9hr3eGZCLFJM3jp
GNWlF5hG20F4JKtwweUPI27OiM5u9Eh23yUVNRNbLGf/A5tcQ0Lvr3wlRZndSaMe
A5SzbmY0dH2ttcc8dh/GiKp9XpEWBSF2lFVpZOZZ6sa+SD8uaGy9oVRP5dM8Dyyk
8W3724tdbM4Ly5SVoSm8XVhiQOXMyPVj6Y8fbhADTuVMsGO4xba55HLAZIb7F+LD
xSmrKp7oTWyrtm/5t0ckv85c8Xtexg4r7QlqNg+6J6/Se3In9B2miuZKCbjb59M1
aeE4rjJDghbikOy1cRXQCVHw1QlBSbbXRxVakVLmJVpzrOnGUse7X3IbMEsZKA93
xYBsFx8ZADjVG4q7SbsCmz6+li/z+Ja0vz8DzEGtqOPk091zGcQr3atfRdguSBWo
ZpEWo3RC72D8inzOHwVBl+dInIQlsrdLWCi3Q8ZDQuHmIhNpDs7cFIZQd+2V0Tel
iMb3s+SgXhYNmjmGxOAcYI0hbUL0kd91uhND0isNM+WHxmOQgUS/NOdLKeaYQrKH
BYxwpa/Lu2PDOkffArOFeshYUMYdav8J4Osz06rRrm1Qw0vKXkQbhQ2ZLFLLgp/w
e8JwOndfOmMpsD4Q3Cd3u8EqPWVJtxTXUDjPYq9rUBf8dqmVq1/Y4ikpUvNPrJIq
lGTt5HAZUG3ozHTz+/Xds1gTtlV+DmPDlRTeRXesURa5UGNlENPeGC3tBLKbCDm4
6jJ5+vKMHIpP5GYfUHdqoVJv0yqj4iAhx2LGBjlVPG5LlmeH3OuDBi1KXKMdqZ0/
NZ3WQ9WaUFnzf9JbqWpdNXgvWjjBlevs7m2MvrWF5NQeXGlPsrglvhqsn6W0zeop
76VIVz1UUi9M4g4msbUo3/IF2eZLDdD3z9OrJR3IanRzSzds+gIxgrxAh3UFv6XD
8M1pPJ6sa0TbQ5Ki4zkYrWgfF7Poek+StMiwL9Wu/dFjHDgp9JFUS1tzl4Ts0Jwi
0JWDW0ZsphSEosuIRSdTXcpCCeMTf5EgSIEVlAbDtLM5LXB8rtO1QWGaSvG1xQqB
0ZGd/wsb39D1RWAMMsUpZ75fa6AUJXBFaS4GOU5uMAIBjfshx+3uN7Tr3VzMwqE5
DcwG7fAKVrFwK/HE+wN95orN0dKT3rOLvAduZeTw7hcsT28WV5A1ZI+fyBJcU7hW
8DlN6IcqN2C8/+5/F7q6iSh6SK336mQ+gSAhIIi8azz8yo8OECO6avMCfVBchILd
/boctPmZrmAGmYPtBv8rtQbIelY/6KB2QkoO9r+Na1g5v5eufVg6GvyadO1H+yLq
T/5un20PO1gm5izzf7mwRanXTiJqw8v58F3DIyXOpdbjzqf/9IGuxeHBxVyd1sWn
H5lScVAOI4A6e6uYpHL4XvrJcY42hcO9Re8Pa7jQdRTY1wo+TMVCBgTxPcuxg076
t+y47/KY31840ujAZTk8eOJbpzCOMv4WjzsNIGGRztSjGQoWciCHKx1dZUZjZRpK
kHM0mhDMnQgktZC9u/mgQYjRevWFab7rlqliNMiJO0/7ZYBCu6eUR8m28uLfu5lx
/4cuu4q+7gRW0VPgusrq2WZ66hO+Y4w2yewHzDx401bs/yWETMOuUNXmGp/dJVNo
Yy0Jec9ZCsofN9n+gbe2VyRP/1wxGAYu8jZX6bOFwlEf3VD+NeVpCzk8VY7T9ya+
HnfbL4wNOqVNsDITwxbLZb2aVqow8rAQLAgVZrXDjlPHwPhfxtJMM/tpwcRMV6Mx
Mqxi9MT9B2jMJU6tjm9UV2fZYMedNn6prUEpSrP6Qy8m3gpktqKYY6BgRMkpPrzN
iQ+4lpdN6opDJBD6EiKsxulu2J6k0rbmxD1AWJAHbF3C90pXSQXKaBhgcrcG3Opp
XXTuzaqWlujOp6Ovn8nbIk8mKh2pC40ZSvWA9FpnP1RoC+uhutUcKn8NqUJQCOjc
cDKRZyvLdglaTssc5hOjQ9W0BUP/WaWZEncZG25PN4D7W+9cTWuoBudO6F3DNAaR
YZI/aJRRwDXYqwTC5Gd0RSgg1VVMYuRMDgfhoL6Jsv1I2AddxnzGaQyTivIjjx0k
2L1Vj36vy8lZLzP1/XlII/krMsirIJEdDnmWEflJN+DLsS9tx07RJvukGi3RScip
7Izyb4/69aWYDZD1e56ACgxxDSic1lDkYtTgYZFW6B8rUuSmrSHlGcwvkOgXx8gA
VXKaixBGWC4qb0YuhwfZ4KVf5plwAwZ/U2lOgiYqjj6WyspINtrWgtSQfJpEG4WG
ng/yZQe7Z8ND18wTJ53TV9st48vWfrW+iiM3OnkmuxjSTZDYa5+2fc8bquoQcQak
1ozHhLFGqdxm++XeJoNTjSbnE2BxuZ9SHwCsW2/LPv+PnkGlypeHUuf570lIdj46
zZEehO/lvMWr8WyDOFafJ42v5VpegsOb48jiwoZxwymROH3IehDGCptXff5mDgni
aNa5+KlIQni+DF+Uu9ujFzOnvQAu/cruHIVVnWiT2uceS4JQpXSo23a5OkS38xM/
NLo3+7BrzEEOa/J+Dh3ClrButzUNCdhIndKAc9pVmrsL4YFHf8HnbjsfOJSuVyFr
EGnu9SmePhqUcDwS9Rn4didqNcZCzScf1KcShiHmnAViLCGyMhbRW7oR+5OQUjqd
gNTBo7pQjx8RTNS9ZaCFg+hm1pxFQYuL/VisHa3c9niYhYN207yI9njIUzWKXQ4R
JE3IvM9IKH5yrdO/v7WsrsTzp7QSiY4u/TFMF9ADAXbAqHM1XRBkn33+fHjZZUHi
wPbz2S5jEH3WLrQS3KbOg9C3J0QyhJaG21jAKTM9Sw4b1PEp91HjveBxDv7ls2cL
8TvbzKTNiZqai5zqcSGluyXIpblZ7I2ZOGbff//DZV5N20d1c26uREmrI0DJLKLM
IqekEwbEp2oCj9lPBU+r+ZHW4SylWlOhtK4Pb22Vy9K/eeLiOIR3ej+ha7Z9mK7U
piZsOaABsC0GuxImBEL7izxPZGfXN+9KPW80/499mj+TVa/QDFpfrtzbsw3LwIvU
IbgX3z71TAuCh2kAFFhW88gXhjB491L6MKEZajhdR/14MUjaoHdfanqqDqP3V6hD
O7zWLuXvBaFpd3qboT70cRuhou2M+r8+vCvYKlB/TNx7brMxtv5X9zyPJ6iuq8gx
8KLUNzVeP8GaIkQW/qRe86J690nbUALZAWl9aJnTOCqsvjqYyG/LAgLMuyv7dqVc
67I/1VWIS9bz9RTLAGs4vK3GMmEqb02/I/yhXLyCKapFWlXVvy7NV0GKPi7p5yHb
h2ete/Ck5+5HYxcYnLhRO+cctQ8lF1vgyMhTpCMl1oP+fybp0u7bQ/l1uP/nZVDW
CQMo98vT1d134D7CtSU+Uzvb/CbnfSDFVcbBXqWCUX71P35mb3itLU2H3ljvNyP/
eb5Nj3t0Cvx/nB8NzWZcd+rDW1WB6E/2WfsqbHIR+muQweBtRHM3f6BIli9peGwy
T3sJBYGctDut7ewTijr30LzW+LdQZFREVPpAgTGFOmg+7W5J3goZCaFZExUNSChv
kcWJI6za2zbng/RUNw0bxoRM8kw8F6H6n3B3tP3obT4sTlmfKIjJ9a9SvnNNOG7E
X6bRiufXzgmDKCFzrM3g55XkT/ATtI513KFmhZ0+kFG7IZvTUoUDjTG3KUGcLjsR
c9X2BtFxemQ4pAi69rtXIo2HN9UKEYgDM2XldIXMijGk4HIfDjNSaZyTKwmohsCT
+xaLzknBVKy0qS7RsSD9gfwgZrK/MP1vRZQT58ofRoWT8YmHhQe7H+n7zoOu2SY2
pdjZxuHMsZdGrg6L7vdhe5LAhmULMi8tqI1Y3856ju1W00wfA5CPv/CxVwR9Qv3u
Nm6jDY9RHEAhU8bE70vz4khj6Ja16AGrR4gH38/hDB7rUVfjeQWT5GGbXVYNM82D
cZTrDqbAfXVVCUTVBKrzXUgdSTNe7L9LjckB2FTxJG7Zzdgz2Fpzcy0or4DQvL3U
DknTgDC0EpcwfCdIvUgnmSGwgCjC/TGUlprlZiubeNGQ6OvbHrKugnYU15hKy9Na
MUwcDGWsCc5rzp7mxYSIyPZpoNJnZ7aGRa0rMiM+LLCRnFAS7zvdFK/d+/7s6ANm
x5YwNtJMsJaunhhjA6m3uFNpdOKPHKR97BAiZ7Ty/auj4bxDjUypQBZmES9MUQnF
yP511UYRk3AXjtQ1pLfozIqU7urk+9P1kFjtSNPydVSMIyC1vjf/AS3MyOR8Bo5g
cz9BaEwF3iwUC5GnehhSfsLVpN+TWG9E2mW8CeZbXO2TR07kedcH0o1JrR4EIxHz
c6MPK3Ec8ndUePZzG94fMo7Rw+YlyLJ9OWTmbPTiqECWDomA2rcIlGYpKMcuI5Yh
DaLv9gmNX4Tr03i/OZz8+YsHBRrzO4Mh9m2fMDgYT0xBZ/EyQPoHcM0tt1HCRvjO
eB7lfbBHkSSY4VLK5bxTDl5x6C3kF10ThfoCBn488v7Vp7k2tpJY6fuT63r1XCfD
IXOJ2KAqLRnw3TXtVwNurQH+kzBALxVve6QElFW7yRVeqQrZhQkFtvU8wxIzJKf0
RxHPXchX5R+MSs1fGuN0R1w1eeOvcwHByqJE4e4av9nZW4CgBiJkvPPB2ujO8FsE
ndv9zOYAljOnHootZwwkivxGT0mJZA2IxN4ji5y8+XGAi+QnlB4kO08egoKo/2W9
105IeHUshoaEWbybw9rsMqwp02h2D81bIAgB41PaTh+Ceoh5GVRaIslSO4IqVIBR
+LhquBrXV+ps0OMbSYP6b3807MuX3piCIRkNrff9N0LKY/TEsbZC9XSwVCBXQCRF
rfD0BQ2EfqXH0nz62edwg8LmWveaSopEdEf6114u7ams78a2Z3XrfNfjRhweyzSD
00HTrzEK6hrQfgdfY8B16a4Wf6z6kEekPYuxBRFsmUee9BXY6Ag1riedY/qIY8+C
rrR3LO7pDSXMVGDiDd5C3ogt0XWV7eM2jTnaqoXEmkTdviBO0coB3ItKyW1Epopi
QWOP+2b8agZyd6b2etWNuGoO9fpYEPMIU/9Fc62m6TQe6u/6k9UgxGAlKvGv/T1E
Pwfde7xiNuW11XabLOemWnHcuIS2AQq1YMZNj3/IrwOj/1r1tzN+aMYvi1XGhCMM
6P0sh8mjskZC5RbF9jZmcteQEhEVNdJFsjSM5PyEF7sWY6zUzlFXamZ5phbZ5Epl
n7uDk5zTLFk/W0Ifa4cUrho2kujcsbqBIGg214DIW3b8/6Ea6RmP/8hFdp/DkiV1
JxHyPcRFEgcp3vpOb67BvgquKgHeLYY3IPTDcG0+bxX5C7N7nMI5Pkq84WwxzSWv
xN+vxI5P6ACKMu6lBcHHPJKidMNl8I+xmn+IYznNsfJzvyFOchxHO61XUiU5x/2Y
LFqjdUFJ2kENvN9YywJNE226/2yV2r9Ud5dNbr+P5K3N/2UsKnX76pwyPN4hcxWV
msXe6v2zwNd/DjhCc/TgYF82fQDrJsGfJaxqpiRtj4TxvscROSPhPjM5EB4I08fM
ZxzaUoJO8/i9Bu9PtyE426RgqxhkVAwPUAtR6GM/y2O78cGvxk4K7w/lpt+XNlUC
Vi9EBbq/+51FRjqc22Nnvy/7HAJHsCRDlUKy2VR1mbLY3YEXSrcNdU3RM3gQfkem
WnHly7DVB4WfCzn+i0jCGVjCcKQzOLmX4ok0C0Ag4mWNHZfZbzlZO/iHrTeAH2Xh
k3Ytep8quVG4YXZD/SNFNp0VXvndr5AkYdNhaGuUTJOVoJwLCmT0FxUL9TyaJstC
HX2NSdwdGdIMMEolxvZVUhKQ6xzoavlGyQ0bAp3wPC7kYyuFNS+AR0875Ma7BjWm
esOkvWG5MuarY9VH++l3lQ/bGOFhVyjxAO95MHOvuB6Ri88/itsd028Kf4T5Qs4B
2cs2jkXSz0PqgDtdkGIattg5VKr72izNkfDSbnXvM6Rd73BWT5W183PidCCnHi3z
/4X0xVd0jdbCpD2mqsdJT+0QKWJAnP3Xifrf/AsuXQysKcZxsiaADAQwG665XZY5
MpI+vyBfkp5+FSxBkrN/xSixkbnY/CICbR/gWIMUEw9Kq6NBgpK72QuhoZbCuUt0
SHmecUgZHzBsX/AECdbNkjPDryQfr874PlxhB46tnXo9zy2r32L5NhnWF//aLflk
klbjiYb0FwhkKMgRgwi0jfaQrEr/7LDB45qBF/d/7PPL1TWWNV3+Li/2nZkfWX0y
d4pJ7Sci5PaAkVRru+Q/CcTcUAhG2OF0J/Gusxt2gVLdFWuGCrCzW740SWTdezyp
8hsbq7RU8IPWLzAE3d1upp2CKnwL82aY4+2BvO15HsgMOnwtxXD6ZiJnsDHOkEUt
DwAG5dcGA7zRdfBw8YBiFIpt3H1tHcLbITSWy4Ti7xYUUJ1I78xLEsiXgMgdFC2e
XiyhJTMQ4XCVsz9TpFvoDjhvGQJOz3OFD+vS0C0yLgDvMIGJAxbrILbxA6BEPnj/
8cvhYTJSOkOOKZTD8c39W6VZSykkTaE90UVL3jKYzi5ilQDJqJGTU862wZOFt60E
ep7jyBdyX7JRG/INoi7pvDCeb97EsgqaAD57EB7kf5J3vlCVLQghk/ZyVgJ6lCH8
y42zMRveCyR9vEcqoOEPwaybV8pQla+cStySjSLSlkjPTW0lI+txgPpjZgOx4Lgc
2yEeBLoxzGKaJGpBDZkpCXC93HHBB/z2NxuGmfVWwMb/2HHHcy2mMzbzopzfULcc
SV8onyqidn8PcNjQqbcwqSV/tkNxRu6hKgYo1rTFSZOESOXctPdSlMUufn679tUk
iz0YHxWBjYP/2/2eECOnKJAyzgBSsXx/a3LkMKp8zGj2Qhry6VvyFuincJl+K+Cn
ysEkZKBrBvgkbnWA6CLOBL+Cj3Fuk7KGc5SNK7/S9yrbl5jfGk6Jap6bzN6Kk1DU
6NaZ33rkwYEuMiiVQr8ZfdTXThPAGYRGUJrUdMWOC20LKmdj8WkmyFSz3hqah5Hy
s/ciamOqiNSG4qSW/u1AjON4ogqF/86qpxfxIWktVj2fGoSIr9jRLCDjBrwFN+0B
HfqdtKlkkZm5lTvgIqaPwmk6LvRhPRmizTnuyqSDnbDDW5r0zIEjIyRcj0KgIfIR
MbcM/IJkIgzw2PgL5vN+vtLfqvox8JV4NlOhpIdNW73oeaG2Ou8CMiz4u2byJdkw
U0+eddwjpgPdd8MltTdp6Ep0HI/Fu8KGwuBJB/J5XrBmgTHHuAvetIbJSY7dTrHE
Vvchx5iyqwPITK9v3DUiYg+cfJ7ryRn5Ym6am0B8uO0CJ9vfg1R9AhxRazJwSxtx
dGV49fsajNuQRI9zQsY3NK/X89xN2Nykh4t64APUah1+w1rN2gnMPh5ov5qLbzIM
DuCygv9xS12gdaxKBgu1WxqdrIRnlnGjWcBdPn4P53n1TZ4fexr7p8E8tbuLnqJc
xkJjTfYfM7qB1rXdqk9fpvSBVYyisGLR+pImdYxxvL43dhG7oseEkqALvnA1F3Aa
geJB9OGzXRWiFuFaXnMpbJZkwWTdLpvqIAG5zaKW2z8lQ0LfhpAY9a2Wry+74f9J
E1JgHgNNR6WkZa9U7Z1wDaBfH9Nn/mvqJ8P3+nRGUzTlCtFymv3D8qyrz+vMPNI5
j5pJJwP98ZuAaml6Sy0svHCu/zhcXAGvPmDAdyR3kSN7KxygnOcsf3kF6Ceuo8KY
zfTb8mqiKXJCdprcz2Yk390Hih6RgAAV3Z7F2DSLB3Dtiy/Pu8px6wZFgsbVHPl3
8GAoS0wCGlACeeP1z5eu/t7PJzMiWNJxlCAvHOd2Ivb05ucTu4eGoUXaqxbeSnZ1
y9hbXU/5/bPym25chM0WKFNkCXhZsNbY2CM02zKti+e4wJQ3CiBJw2QOHKfBEz0f
8JE6RBu4bU8ZQZFQndvGH3VzuGPjc3RGDS/Kf9dxVANthE1XNozJLOCkmZtY4Kwc
Ej4s8O0za5gU1rGRqEx/xrstztfK/NNWcPyq0Z4agzsSd3yORwv8xf/MgTapy/eO
/V9QxmKIo4b/2wAU5FifUNlV99X9z4CZdkPImzIQxCmLmetTuyxpeNusEeifDygc
p+M1giJAbBpau7BfGJoz1VwggRpixgFC/iB+zeVqNZ/LUKXiNfG3eMuxvvSgVt4w
g+5slL2nFBSOFt0jFrMMHaCmNLHlsj8dkRHC/8Nej4Xs2QmRAonlqV1+t759hGxx
GWGWShO9OyEIremEE7YKAr1hK9jdC+8Vb61ZmUEn+1jnNeDdJIf0BCzZhvvzGDrd
1z1bLhRJXTaqqXhBk6XcpuMUsYM2WtDb5OWvZa02ba4QxReAqkArsm39ZENkpgXq
vn8b5lmWHbK1LGAQY5uHvtx34Ra/rc4vx5aYXxOySDY61l9URqEBwVLbL11bozsp
76lvDPVya4tiKMyGTj0FphrNiwMDyhd4SRqe7FppRCPdRl5MhEolHDbH+NXIDgrm
9CvF5G/LIaeJUuo5vPbZyYJsMU3GC/nuJ2+xemrGgv8sgJPCCWlaEbcYASWyVi6x
J84q6p4JBxZt2Sf6Nwm+wcQ/RQ+7kSA1uQJWb+XfcpMXNeuo0lACpxDVNIeOhzgi
2Air4zGb8Mude97piiyThfDxwaqKZY6ggJLFdT2n4coB+oZzgEzVhDrBwEkl6bT3
2RhY+/D8818l4XL53DKeDXLmiBfyj1KdrB0eV+whNvGqJa1rqpRQBSwBhwB8jBB1
uCgt173crqZhr5Sj9oxcmvyR6YkwkpzHIeF5g+pdfvVjfu6BtHKsTj01ZHRT4hWh
/30vzjikU8rDJIqkwO3pynk7hNlNN0UK4K6p2c8fUQo1l/dNKafloig13IC37i8v
huvKY96a6PDDXCBVl0zJxQcFus7v6WUeKPc2epjfsyBr2+4/2ECnR6Hg4TiLyC1L
uY3F10XSmnLpvVtErYFwLXHtImWMqKSUBcdqkn2dCfxbROPYTBEYUaGSFi0cyH3l
y576p4mEt6vQG5Z6RtK7dqLjgm62cQJnRoSNV5OeZXiMEaWt2G5fAdJoDjiPIy7Y
gWizSNpVqOLa7J87BUq/LSqtiQH7tirc66gKM2/3ooX0uq3VJcaPxK8Ny3KIsBuu
MQaTS56lo0JXVblI/2r1ngaT7wbOT0Sl5r1+oR7NkERtg+N3SawQFSneJgnpU8r6
2qRxPWVYWmIjUxKHATJFXRhpHPLzS3jdEoJtpGAClpQgr2np+/N7m2zon+jXg5EV
xv+tYpow0rEVHn3ZR2FIAVD0FtcfJgyEhk2K8dmDk11/JLiqAHAs+HGHSX6YO4m7
prUp06nKXWeC5musogjevzjf44MyEyg73WQ+HVDnwe0tyqdk5LKMujig0IsjfAF4
fc7mvo9L7mxqaKpEjUotewOJf7m0exRzVWJej/BiMQZUUS6m+F6wkDToaKtHtUL8
M5g71JCMjVn50NcH5bftUuug4ddWEIGxs7k0dAh6NjQTkR87jt9W7uel5VWxXBLh
tFQPNEkPdJJB4APBnShmyqwljb8gTSe1iG+IbAVD7453dKa5ZePjbHprrU7ePg/V
iXrEWPJNaIEr+TxJU29nBdsEXEbvSCJhnWpVUZx+YpgezV3nMzKthKhzxN+Hc1pe
Fwb7hf1ZGLokY4YEqq8P2fzS6GCi5MlA01sYRG5Bh2rIkIaFQhUG0//oUFLLJ/7q
+CbSafBbPk+quP8i1NQ6/d/Bt6EMRHlP1cbQoFMbEhLHlBVqTc7WJHfTwX2UwuU4
RCNmvQfusZ94NTwydnsXayCi+Q3g5Ake7g0qi+62dcbEKOhe4gC/sEabO3J46lA5
hds9NSaOVfC83u6hR3Udo+1l0EWWDnDCezNYhmWk0/+DVsc4krsXE8Wr8L4W3usM
uKjFxI1Vb89IRJMYoJLh9XMqUhWwW9qLCZX9+6513lDNG+lrbFgKd4B2kYtChHPj
j2HGL6OyUTD0P/OviIAQNpk2KqJBNU9UBjmuiIwL5eFDnFqicYK0O3bCgbHF3Rz7
vfjnEuq25/9g3L722PKPEGEbgb75EMpDiKty4s5ngzsxfIhymeax5s+H69O/NLSe
dMmrUbdzpZfz2j3wc9NP5ErMNnWj3AnRQJENy0GdDoBeEa5OaMTL27iuC3ZfxEb1
FQA4Xl8PsI0STsyXHEMJZ13UGgCh6IDLyrm6lL+owLzQefySUNa9DPKZZR4FsCgP
7gSQaGRDbWaz4hNLmiOMB7VWV1lSJBLii6N6mn1vQpQHWyjViwVJs31i4ySrh/hi
oAq3smBmsptHbQ8+k40Fyp9jjQfKRPlMdy+RVB1IV6GZMo+7HDXoH/RUD1CCegDy
fY50K0vsAFcU2j+nTJ1bIm5noz0UmEUCdp0T1Z/psr/fn0/04ug2clBDKJstA5ho
m2yA64sg4c2WhiMrXg+IRVqIkf4jmvKFYoNfEQ8jJ4e+AmMuhV3FXu76xi3WItCO
CuFUxaBvPBwWFfs9cC3Lj0a6IiHHRYmjqlIvp/8wrNlJUM+tku4lp7xztUqzKYSb
6ZAnRzFMXhy7Lo78Xgj9VdTuZDYx5+uXl57/Q+c28EqA1RyPJsjHlQ+XGLhFYTt+
HNvZFBY2x8QzcYUIBhDNf7ljgkz/56OLQCZ4dk96+3aX9YLWpi0q6dbvvs0mYyhb
NPy6rFeYa7Yf++nXqx97lB6kv3DD4VYK/UjQUN1XgdNdxomOVOXj1qcI9UPcS4ug
Rjb/j/7gKRPx4cxs72oqypMSc2v3ItCsmnCtds9ijI95s5QgjMmwsRTEWKtXazn1
oCHvzxb4COuJ4m1WOSDmqQj+Yu7nWbJpepbwo+0t2lgp0ZsHyGBl8vQJJanhKXus
h2aXhIJPD6vSl6imkcnj6BKSg2ri/uB4PkxgEe7kkPTQqjyPb5y0gUkrJqrL0HAL
V6zpHmWUKGU818t6jXakDVohTwYupW0plNT1V+B7YN1fZ2L4/gYeT/uNg9cjewNN
D8w++zw8C+FXP43aT3r21UXbwspv/l1beyhxIV6FdYhtZ2RhXyfk7iP1Ldh9nLGo
GZ5Xv26QFh3pZ+Qox56vrxNEQGHQ8SiV01ci0BW0Bbh0jj727sW7aJT1GkhEj44Q
0T7Y6m5t+7qZSvlTBbrrlavfVwR8DGsIHHePkStt8h8XR+sxKX3vzMkMveHYnQmy
B9x0NQ3IzC9U5D7r0ydBY5c+i8i1BidjKblKrNYn086cL2Rg63pwNIJPiVmak3q1
VcMV0aci0SqwsUYKcSxrKJLWThGFvCSDN0Sy4Qokd2BgSP4Pb2KNlp1nQZUVmEiF
u/tb7QURyy/OH9Pu3+WpWjXFj1eDXi3yjhgmd2h6l/damSll8YnqfCfgP5kXdfla
EEGhUInl3wtVf5FwzSWigKzFJlzMZ7EGhDjNDg1I3vxWFQBlD30eUE8Bz+hZzIxS
cMl5tZl7Da1St07b8TzDf8Xy/KQIROpveEWxoJ92dL8dDdveyhQnM9SFHVPhVcyn
b0p3VmA8pOY2Gvg4Vht3+ZA2RJbFUp++mnqX0Z3eXb4vKJSjGm8bILfnCbD5E2lN
AwQdH9jeYMnvQcT3eqFiV/k/+N/xv3WUkSTJCEqzKdButMf36ZXMeKYDX10bEAWJ
uCFytHM5yCGgMLdy5nQl3+lPCRDnRf/h/So0Q29XE1WxQYokr9AppVjpWrRIc9Be
CrSKItk/RwuAtCtVB6ztq0L/7OQLdB02BcYtd6uKXL8hdHY8ZmYzwGz7Iyf4Ejgo
XoAr28BESjeus26lOhtKJAEttHY5GPqPGP25pIAs9+ypPCe6tvzPMPdfWFKo/atE
yCQK4gqzh01Sc/XkzWvLe3vbbmbQ3FsykYyWNRnREJ006tB+mwGqRKkcg5V+bkTF
DWgiTsVcl1dIpctBILLTx7Fa0V8IN4qHdOknoSBkaqdsHsj5+sLNpZ3guj9Hvlj4
R033fiXTv/J0TwhvP7jYw3znjmrKfHkFE1ccOBitKmxtUyPOuU982bWDhKu5zXHV
m8Dg9uE2YsL2c2aEFsZgN9y4/IJ8C9PYuLIFsHAzHcMbyk5EEQUj43UlguvqrRd/
AVVPr7TRUkBpuriOms3BDuFJHOj/scHUxwldOnrngFuxsQDHUUAVF69tGTKbHTrx
27lktVhi06Vr9GhtvoaGBbydYg3pzasHqUNeqo2zor1jn1sl3j/XQJ/yCpRpelsc
6YqWuQgE8bHt8kqL6f68UznIG5KrzBFhQQazgJFHC5snQLqGbDoImylAKqhgik91
8B1Ez/WLyFwE84Xirby9xY3aMbAUpotNBNTAkRn1GQMo/8GtakjxR3qMlQIU8nZV
NF3fbqcmEKIZu69KSZmYVeDhrKdtK/9h1dqv3TgU9kfCWlrvAEHVNtjb/jHHJZ+u
to+ed8aGx0ASusBY7PfzybXAubQj8FmSjVm5GqIm7s3Yx40dsXVMpGSkZddqBAeW
t1SLkIzRy1Q2AVCAE5baFMVntl22yIH/x19oyCx/nVCGSBxkTGhTO4kp9eFZ0vMy
kSMejxTe18qkeGlMbh7rdpJNatQ322rDtSKE/Xifuz06eU28tmFoZ/Ir7Z+EmXGU
0lyhH1Zb05oiVi/i/WjNQBoHNiOrNtV6qNadMTnki9UrG9Yjxo7cUiohFShh3GFl
zf5X9vs+fhj3zr4rekAOcYVpC8XZGtvgx6eL3Pti0lHhyrNGC3K1QryC0kH7QFph
dwcz7YCCOGp7v2eySOqv7idIierbStSwHJ3fHdo1zXMEZK6/ERYZOiDv9L48uXUn
+hEx4AWIsLHtddEfXRGVm2emUZJCxZIBhFg8jF1NZAYtt/RFnz1I5kjeQ6WZQqHe
ShMs79y16TrAS/QBypTuedUJho2UMRARcl6pmMdnrEvMgbDGux+IkVNVuMBCmRz3
OBu3Idf8lOgEzXGmicjTgvCBQl12RU9N/JNzoCi/GZZqJk0OxWfXlJ60YYeolkyv
3/Uw5EZmDEcxt8vUFhCQP/SaYQdlhcxNNC++H56QannIW6hzGJQdw9s3j2YjcKyX
9TUs150h6SqaHXe6qrTl4ytwmiImS0oP9XEztc4joB8NPQryKT5P3Rwtr3CjV17T
yzfMIGQs5ImJRq/5sO/wsHbyJpdMc+Zfjg8PYpBVyyZuFX3UN4Mb/z6+RT8c3SSv
XpYaT27TJ3lauHyernqx6nHjcLolEE4wKVHFZzLwLh8M3ihYflz1nQzT5tEmZGTz
LeFg5xdrbpsxrPjMQX1WWpBnDIFYP/DYbtVXmAGfhomdGLHNVM3S09tyZ8gGQgvm
CYoMbO0ObyxIdkj2wMJPyIasnm9gY/B/6g5YWB67lEv6Zwca3npp5XjOEfMlo8Wg
Yhvgnj2WB6HIkhG5wwDe9EiYUzP2yeti6Vs6KDu2+5Hnk5drRP9fRGm/HuKFSu1y
BXFVDfga46HBNgQFWLH/16i3IT91ZwXJ0f38k8bOPBNzz7I30AwgH9JHOa7wffPv
gxlI7P7qopbEGTXRDCiRbDXRSxf1t/5yArsC+e/cDb7rI3ORjFabUa87+5tsss1Q
Ej4egIxmBoGWjP6ZMkKwZuS+66Cg2y2cgikbkQO6H+pmXGzYYynqzT/NBOv8NWsS
Y/EjfcZlAo63Z/c+IFAwVOpN6SzZJ3ugGyMPWi86qcheVHVdqVuUDgZJSuevusR/
hD9QZdXokoSYUTFoGuvat3NxHou066dChdXPY6UQlh3eYgHzxLHAjYPoEHOSWOMT
eISu7LKCNzjHK1jPvvKzOsMPXO4elvlU8QS7FKpo0JI2y/BEK030MeNwK6V7yP/c
syT8p1qRDZmIxxI6OnPaFLe9ZLNN2PS72PITy01RVvw58hwm/HNxL1qL9nmwOM1Q
fRr16C2FzNBf6W+kDIn/QFig5EFN/D/yYFxxV2uYlIAJY/O+yhvjBLzGW2+rbAw1
IBQ4jIxpvuhHT6G6SuDZBuHLx7J6dY/49yX8FxlxENXR97SWJYmkMXi7KSoTjhBK
eUTpQnzHgmC+UumpaC2uRpujZcOYZJXzqXSwzcm62WL++e4UmFuzbpRdB11aakMa
vxXX02fHvg2XGtEyOwORvJFI46/YuNtMvql7agDMkXO7yJsKk6NRx4H9crl1nK59
qX/4u/wfVGPtb3EWUjyLjbmqMrvnmBRC3LcINZdetKwWhf/UxNZT5StCC3GmXF+G
vFw4yEfjhELndbx59fPE+ne1IgZkGo0cHZzccl8j0B+mhgujW8P30fNo8eCjmAD+
1Zm/IDNoOGlOMwI0gvGSsNFzr/jmUuCwp44LtU4dGOtJd6QetZNcpuDvCMOPifNe
pIH039oAdkvdOBxs8ar7AkgaCmMKhtKQGmRHwfEA1rcJthNz/RNIZ8Yj/xQRS2Sm
5HBdqddceRz+wX+g9Wn2TtLCe54DwWE5wHWv/tzIow+fOV3layhv9T00LvLaOL6e
FlPX/IORDxdIdA773XR0iUuBbMyVrQZbdjAvXFH6IFcnXr7xjBBjq2qzQhVvLmYV
MUHdr1EhiZr+QnSqECbVlzPV9hy018GXL2j/DeLjx8WpQEbWZvyZYYiFyWYemBGD
xOmTu6uerFGu8rcW1lhmjRp41W3qh+Ryp2cc9RHxVoFPj2j1uCPhFzfNHaYTYtRN
hudgNYdTQxtgKQtMCiyUx8FaAmL45gqwOlCfVJ3tHvIU4nmsjVq1mVe4yvsQDcKm
JDoz4PhLCkbkKnOWAdvHB/7gquuEB1Op0mK2id8F6EICtPaAF8vQN1tbVjRy/3W9
kXT6W3nu+XcxtdR4TqjVWZEzof5icAijfd0meziXesUyAGQzb7IoR1Ep+/3vbJmp
F3Gy94njbq7v1rw+pD4BXzqNn21WKCThVxPFAh2J3uNhZWbBCq/KXhO9swx9YsWe
EvRcuk/KXsx8i/hOx+HXR6//t0fiw8RuteVlsaUIMKcidFCzpdOC5NkGxrD8XMjw
wazHJVmdTAHGUSjH7eP0u/JTnCHe9V7bYltX2M/oEw4EIJB0i/IssvgKzR7XULA7
zbHHlK8xGZxtmakHFRpwIM1hXidhquyJrQdSkPwVLbWQxTLBIQgY6zwJQ5k+2g2+
wiEymFk2KWGdaCUZSezEF2JEVFRf8mKVhSc7Vyt13FbUeKsePcTwlJz5qXc6+3Jp
jScH+xyPXEG5nhCKu/dp2V9JxwK5S6scaNEYXtyLmmfCB3vBh0euw0WKlGplwdur
O0j0oNTnapXlo7PYaWYMw1U74TGMqTgRrsJhtEQrPKKRBY3gqhp7VTMM91lDAbdo
YBsXnwZsL6x7xdfbYzliQtT5vxyjxJXwOX5We9+iwKcNwq/5aH6Gu3Tpr+IvvyQJ
6PxxWf8fRzw8j9oY7YuWkEFAD/SnssO27tPaziKlubPENE407815pKACChEaEFWj
caVRb3ZsNsYhYHHYtHZGzZWmkIv7fRpr/J+pZpw6trPOP5+36WaT62dn8YTpDVYN
AOQx9FoNkJolichlirO4fmwXQSz5ZyDfjGzumpkIx4lSvl1hL5yZtpKxnNi8B0GV
JCFeoOffbwkS2ncegMb3oSLTTDp2VoWeb4l8iR8eDA5biDgRFZiovf+1AwrI3S08
rN49B5e7Guc48Y4JyrUaTHsXfddTK+0CVvmj9IG9KKw7AJx4IBArDFje2Syn7AxH
`protect END_PROTECTED
