`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAaLTYCbzwMa5T+vMkoyektXKcw9xb0mY10yURdRIDRNR
iFoC3tW82Q6WVqC6B0Ta2gG2lBid+9x1fQgoZk1VM9ULziVqP48CduAyi/eloLmQ
l/xysnmDoeu10EODBAXd4n0fViAIWz1Xgw4yX5S55d5f0tbF1vUnzjSJ0Whi7yj/
PzT8d5TNIwd2f7iUbDbgZ1TSC3Kseyu8JRJ4lMbdzTBTBW+pl56dmfLSLTCzXJHa
19cpPwTyRQElErYb5oCGplNS7VWJMKJZ10Ius1+kVBZXzqJ2J2XSSO0OkLdPNldJ
WAsAepunNr1RAPpd3M/SvTAavNL/6RDBRFm6iN22sgIc6fj3J+bu0iRPqOE1T2qv
OURFsXtRZOtBObJEjs4znc0AITVE3uKEhzQSISdH9drqRkVYYLv8qhN2N8JiZkZe
2gnYUDRpPWVwB/Hjc/0f7+VtNNWOehVqwzcZj54pex8HOZwQJjrg9N/j1DTOUH/O
OGeLrF7k+/r6E6t9q0I+haiTxHBq81WOyi08O87FmovIHSUMvW+ywM9S2mAB45dV
CBhjWoz+vkXIwu3qSRbjnYkkGHe1YIDMYVzaJihSUO0+HO7WU9UIQyvzcoMUOIN3
jvFTt3HtqvwP1fxVZvc9uigMDXAeyns/7/imV2CyBpkNvJFORkfHjV8kbEYUxpZA
MmNfsWFH4mxm6+TIvSb9CNj/WqMeeBWrR4CX/B01vo+hTxJEYjC3EMw6o/e2T3ju
blH+gdmGma93QZDhDjyW2aHVGm7FVqqkpUDJnLdmQPfErzOi9NJgsPZX33KAFGQV
4Niazma7mQhjr+jtXhxtIBv8EF3nmmXEnrdTPsb8gugqZGiXcplUlyTR7ir8rSE+
/iwUH7LxCOkVT31M9R3SxcxyerFXbqWAdV7etdInolXSmfMRoobKMHCu0dScxmMX
0DrXZJ93nn4ypIgktztrlrNAurbyoV1fp4FrycWkHxuCiNNrBA6/cYmtK+QMhTcZ
3PHS/ABAcOJPUP3gaN+z+F5wD5A3q9E/jsrZB1SsnWt3HRFYPSW6lj4l8+cl6xdF
5HqZjMGQQrw63N1euJ9Rzp9guby8kiuYVfgbwCa+FPCwa9KznBa9WdNdUjTJudPH
vFd8RjEKoQJTxmuS7kyTyyOCdhpxXLWwo91rrgHvFxJeE9/Dsh0TmVQmpOUyridq
ZlhAV3AXQk5gLlagfT+Mv1L+ruYMtQ3MRmWo8sAWKua32g+jFzgf+V1HemErJvcR
X3y8CnnltvI61ywp93SzY37ZL31EcpdHhLDiyJRoB6bNGe4Fr4UxNCgI5XNcuXoa
OuDNOop6CzlYNSB/zOEYlKYPoyf6R/tUMuLbRuNwDS5YLh7ux4UBHkbw/RdltNbE
IOpHlQpvT6idhcibtwQQWItt7kWTGCPy23KAcY05ElAoTabZos4+fuBZFPNTOxMd
puvEGWoGCPxDO87xtVl0zANkPI7xlUWRDYShxihP2kmDUi4J6DUnRgKeP13Y6BK7
lOvB4Bt7mgrwy+8OtdojfKFnBJ2WXzhcxewDX9rYYEVfBoIyWuEs2pnPAn4FW8SC
e51CRvevG1yfqO3cuvMHsOURETfwwVyTssMDYH5D+KF07UPDdoqLxqyLHdrEm8K2
xfFHPnPWo2pMAWv/FWij98Fx4GtW6gZ6th+xDStu6IcgAQC42C3+dd5yXq8mlGcy
RTmylgk7U49bhvzAswfDe3MyLGtlN2ao9rgfUBJBI4QrI5dGGSncbwqJ9JPwSm3F
EYHuoBNaIcLxXS9KqPMhBztWH3wvPuW/OSuOWKQB8ejGR7/qxZRUEiKCRYUc937s
iRdqcPtpVPv3xQuXCCFzAGrGIuBciYOW8GbFN6dlCGzK/SvlxiSLiGy18y8Vxi80
3pLMug8DXulHLQNWLL/sOFdnVtH49NeGvq2avBa9akingnq2FngksH+HZVF4hsjH
wrk5L3Outjwu3xEy+05CpflGSD2qa83/SrVgt2Ts/quNDcSzRm7VkIXl4e17IiWU
f+PbXcOvf1+B24YFVljdsRvpAQkp7vx+XEoe89gxwYP93QiXCDVvqYrKnQLIdoWQ
vzCdZDg7EBXaXkmzX1SCSblfeYXNvITbBq4EziXXnWilYUi3MVbHsFFRHOHvhLkp
Ay4jiyEbuVwC+vxjMeQQYMj7+r783S5CH4ClCzTnbnuoQU25253oABZ4m1eArVwO
u/540dAwAMk6gckZBWnTjbgvNOao5h2IYfZkkcsc/1ivEgu7b1fhQ8CiPwlTS972
apIKezGiLE8KKYxaFVpx4Gk+c0haGRqulMISoYHxyAnJLY0FM+flUAgCU6yMDqKN
6CG21OcFmrWICwNBq2S6E6dKYdi9Cj+7c/evawd8uRulqOXYkVgL71p2KrhasLpX
bC7rAwYxOA3BspcWkYoRVgOaa/wxQuuVQ/pSLvPBbu+pbc2jOo+CAoze4tEt6ER7
FVtZjf2un/BvKqeEV0wlhVCrdwPGs47DxGmrROsPUpZiHWlGToxd33XLpkvfenEZ
JvnqmXWTfJy+ak1oHIIzhuCA33dOuBMEc5taxQFt6xPbtyhrFiN4kYVOikMKhM7z
1pmF9Le+oS8G5PaOH5VXPsJnMqXPskHY31aE+czCU9Rs48Ahya3fZm8dMYGZdtQH
dh/i2noOWdfDgEpGDeyZjEY5sweu4dFRVERhDjPpZFzc4bk2jNUFmeTv94hYIh83
JYSIHpn8UV2YmD5xQgWU9HeVeJO8CTXQyxHYrhLw7qAoNoWoXTZL8FgpijF5R+bV
l3WhmMRjBLTkTUVAyp/PG1KNkreXM7CQvrOhKfQdgN35WL1ZGgk4xbSYX/eSlEdc
Kr/5pmTdgzui7ibuJLnZv/p8k4GFafc8YFA9I0jAd2jf3ckVFKPmvqclPpGznba/
sSr0o37G4likXjBQA0M8LE+gHZ/dUkoRHgjeVH3YXdxXRM+o4ckkX8z+SOUNdpU5
Nph9zEHVqO6G/+7ChJqo8dz2bIMRXqbnkk/GaflJE38RH2gP0pr0q7RjGq98MOWb
aMNIfCNvTZXzO5M/XNkp4twNO0u7A9/GoyHmUweTxTBQ7UZ0nh26SvzYILQwi3Qv
T//d1siTqzaqoFx1v41lnEaxuhpX0Q8FoL9QEGxFf0xvpiDJ22FeeAHkfWC4Qqap
Zpfgb+awj0mlY2GP4hyRy4Ki0/1Tm+s8D4SR7isxJ1rHJGG4cZ4QM9T8mxaPiWMr
CPSdnRYoBiwifr202ZlCe4f7yDA6lmDBZeU+3wb+gz2DosBwAlh2GKVLpg+XViN6
p8DMHSX0VISUtK4jqzhOL2xrCN22qMbTRlfgUBKu8n/RRjK/C5UZNKTd2VnMuOzb
v9MC8qj4JaQ7OSbCKxNte0OIT/4wcfsZcaTLrcZojuQd04MAzCLNRIxDVZUshpE6
rnebhp3Wm9Ftpv/ajChG7Ht2N8hHsfRnUA+kSqraX5wEwuZhidmnw3TlA7iUlQwH
TcyF0SycwFcPbEOfJjI3WpbAmYJ/3C86GFItL686w9Rx7nVkXl0UJCEjUuaUwn6n
woEq0EW0FN9ChpPKewYQpwf2HvyZ98x638+e4MB5uPhWELlZxXLE6e6Em3hkFsXa
BB3gi/zFYYVlAixmuv5Dr8ixzbAU586B+L6sdJK+j8CBPct0x2uD6z4JRWJnX7fR
XccuVu35Y9UGGBdsV5912ghyxie2T1EDMCBqwGhGcbQ4tygYdKE9jeHApZ6cbjvy
OioAFVmNuY935ibmCw9lrrn+lfO3AyPVV12p4nKBpPS+fhweDvXCr9z6u9fHYtaT
A6dEm5uWpA1FdwOXqjhKemjS3cHtyD/VKcmhq63Q8NAog3+FeFhyHZMh0SXGWBbP
wtxtPqJAV47b/69RENRz5vAFpfqLdF61wWfK2xiC9L8kWsoQyVDnSnJyiKIXNywa
WNf7tEfRTdeL05UfJEIS9rB4qmaN92WAkNR0WvRMuJs7A0xaC+P3RPFK+hdqiR2r
KQdWd5skLmcrAm2PggH/b3tZE9y/zVSqnyuEbSmSA2EbwrExhhv9OCpdVkwEmFKH
WN9xhMNo1gnL1uBXgd5oeiObuUMz1GgN59dcpZvj1BEjJsvO2vAXGCVEqf0UDmjZ
utTcaBqSUujBTxkbO75ookCV1kOL4JlUyAIpGxKHO7PWsnOM2Mnv6/KYpu6hH5DH
yqzJgvKKhver9M0yD4HnZ/0ktswl2tM5PO1gMVLzcJcp2016pU8C5hI/Y9hh62VD
H1LpsxgpVXvqvJ+m3nHgPsUgA5O0NbILMJKr2I+CSGeDcOF9XFPHoMN9N3uWlIhQ
8NvlL0t/EzVzuQ5SICJqqfRotRA2GLnP7fCKC9vN/kZbJuKk7J302bFb+X7BEaCq
`protect END_PROTECTED
