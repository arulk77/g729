`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
01Z55phGGe5dP07d+5RFWtqrc/9Nqd+eumHrd5O6xfIgAKmkkyZVzPzhUw5ekbLa
rzW43/KntHa7GN6ceGL/MTX2wmoqQGIE8Cv1sdzuF5rtmsNh/ghCAgU6Jgdscvvx
A8Ax+FsWURz7eP4qUIuH8XfQw6tLZ6SGbBLgKAhbAWPJq2AsIC0FJLXAX7nkj3tX
q6HzIbyIHvp1Zzv4x9DVGyiXhyfBkGy0EWpmb/ML4y3aenfZQpXUH52aNTZ8Qiq1
rKeUVrdWn4TmkOpQsN53FxNmiu2omVeE0Vk02qXGuG9S9qC0DdU+6XEE5NwbtiDt
GIAG8AKE0Nq2+Y0TcLAw2+VF9bytxEo4usFTp6xRGy42uIUTOyBLDOR9jT1diURs
syszG5+LopAcKflJlqwszwDN4X1zBeUsx6/H9lNK+R/ALTyl3WlG66vVbZfHNzBU
g6OqlsPNqROpIppdYyNVbIcfvWlJZz00IoeNql7495KblvSU6ts/11QjkkUm6QaR
s2qfcLo58boNuzQbn0Gyow==
`protect END_PROTECTED
