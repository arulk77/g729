`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG9tYhvyZtILvSAv7qrpNUZWOvBkKijPvzGT5XHf4+QZ
9okKvk+IM6cftgcbhYU8WM9AmJ9HfsLDOm2CwyfPEmvtDPuf2yZliZ7tXKX2KSm4
q+c+eSdPZfUvt3FMEybUpXibUjysLR6ODw1nRmr2hB2j3zq8HwssA1daK65P811V
YA4GBUznBZ9YYPXnEu67QTBQdUfkyd3WNnPwwc+If5POdpYEZi9PeG1GCuDnFgiI
fOaSZnEKFanarPJXv/8n1W6lJIfrbiydBA6vKn8h9kajy0s9ZNlnOrx34nSnUwV5
hHIbRu0teHRh8rh5fAtu6+l70hrhojMREAgYd4kW6ek5zDIc/EDWtlVZdc6lUwW5
/kVXdXB/FY8kNoz/b3rVzQ==
`protect END_PROTECTED
