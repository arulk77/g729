`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+BWhzRHwqqpIkCmLv4MOOXYKfPocCctwgzABUtSMagvYtM5haW/mp0gsVPO8oosB
mSo7QPZbOeiQcCrKd3CJxilMBgiKmcTUVksEYFQx9mxqRv2/Nmt4tIAPnyueHBO9
fsUhppWHWEl51nyka/f70ACPViR818szrzbgzea1brtfBShmYK2DjC0QgsG2PlBq
FhQJfPwR6pZQzlot7cP6ZI+Aoi+s+OeHjjiYKhMARtoOmH8rSQAzMTESjdU2fAAG
HkuVrV69L5HtQhFjUQKobQcqmaiPdAoMxMBIJu18n7DXr/g9SE7u0rbo14p/pmIj
UV6m7hoQ7gCO01v5CqYK8D6N6t5A/DyQpNG3fEK+vyQ=
`protect END_PROTECTED
