`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41ZV2mNGlq//B5cNDcl/gg3uMWm460Ino7g7vsBtvK+W
PPKuaNSNHuwS4ZzAiJa6L1k8EFnMkTvFJF/D6m2bDnvK1jiPPMowWF/fZSEnEQoo
6UVY//pyhyJaDCb4k9ZMOCEW6qC4F70Hglp4jCJkq/XK8FWn+/8RGF3q9weuaKfw
dE8L5b+U52nJ11+93f8FI5ULziU22Vt/yPKAPAaMyHZozLYG2zpu1y/FoWUqtG3u
X4VwezyDsN/FW75TBaUAQQ4RAZ5S6aENbympJvK7fSlslOhD9Qy2V6aKv0LaTxPS
sInfW/8p0bCGDN5vSx5BblGHQ+R7P+xaW8bqAhBChfTuGlZm1++1yR9znv0r6T4q
ZaPmOjbWOTyb2M2PCwNF+g==
`protect END_PROTECTED
