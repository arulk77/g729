`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/2kcv1hOAl0zzUmDTnbuublzJPwZAu9h4U3hixKe7g5IUWz4Tvm7xZQK9vHqdD9K
uDOpK2aLqzh4Vt/rxM1JgZEau+31kMvU1KjT1QVcOlLigji04ZMA5g0qVx8g921a
pn4ei/sa/zzS6fl2H99poCmTps5f8LtHzJ5DPhO2ouv83WVwwLYQp43q6fBT/Pj5
5di+vSls9yD89ECmxuPDWOfixaSK1GleVlYAxtmDCJ37JRKWxi1aqyRdJCoDUPeR
ZAbZ/pO8J8BC+Xe3jm9YZJvKoFvFsKampSBDvubfUu0pQxC2kPwxr8PNZ2vftVpy
TcSJCZEi7ebWuNLQFQi4nBiWbuMkK7swqbhjdT588QK3shlfimQjjfnWch+MRCFJ
C7nBfNI5larwKn8EzsulhcOTYNi85E8NYhWQSvgrGsA=
`protect END_PROTECTED
