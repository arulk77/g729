`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAhmeAZ6Tbk9ZtkqFFdlRog1fXU25fE6pkHVEgGpRwRt
gTpXBvkm2V5U/veFhk/7kcqqs59ZHWNfLopJqF6FiqzuzG0erEmR4yQwPR2Y1Vfb
kKJQU5ir9RZwGPhoiUwVQebO3vaUYqwxEDizOBpFgUctlL8hnbeJlw3GQ2FFyqyY
LYXrpAru7PUc3pQSRdcWEVfGE9VPi0AsU1k9BfBZd8A+MeyKYyOHlvm+RcdI+Z4E
5gra1xamXOvkuytMqz/SxQtm6lPeGVlWlUh8Ez7vtnEa6VYvnHUiQIGoBQGdiZMV
1cL1x/7fNRqyjlAaMYGeQa9nE7xE3BCQRLB9PluRedCtbdvYFw9xlzjyz2wx6diz
b12aIDkNXlktxUxbo3AuDFWB9DvumzyCG6O2TdWtBEUdQ27qpkMKfWIFouHWXZAQ
vZ2O/WqTjYvxl55dAdqmeqvR7xJKR/Sz+Qozpe0umAlXjgKtI3KI+ajCTIFWHBk6
1+6D9N8PMa0tqTUqF+/O66kBBM1qzQMDElPtwsH6ckzImIJzdDGf0obDUqZ42VAb
`protect END_PROTECTED
