`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAEWWfdYra8HoCXVh83mbbGMLr2Vnc6FsKNCVV9hNFDp
aoxyjZYxFKsLSjyKLwp6CIRvtvkxAZoPiClnrgovMLnVmMBGLtq8+9qDOZP6qOo3
iW8AAfXyQphapqj9j/+icosQhpXHpYlYTl77Q3aTtuadxsziiv1oOz0FOI+W1ol4
yKvSocdqTH7pkDfBN1360fLSNQjHiu9h/nugJBl002qEsrMkGJBvNZbc54RNMSWC
YnyLMMSTSB9azIO/3JIBPQ==
`protect END_PROTECTED
