`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNOlesGhJP6yKPw2Di5lL6I6RDcKNBHQb7fYuFvDOL5i
lvDaBd8YhxfkblVrHYm5SDgFlpi7hucd+L2gc2bC/5tSyGqZOVdcZ+cdlx86DT48
qk7NTNUwldid5cYBu9aigfpRgW8CTwo+/uN8wP+LwuHjEQ9G0P3zKUT0nxdE1tPl
CU8vNJPbe5iOTLSrfkWcQ0Oow3uASkBaWHsrfZtK4ra/NNE1qdTfP571kooNEU5l
ZUD2KjwTN6W/uSUNhM6OkOMG8FuI5a9T3Yhz4HAFKByf3vXvDnjEQg87OE9Mzaz1
1gUGodRO2rmaZOMf3Xbfp9NcqNsl9oZCGV0jtCqas52Kmhf3sWEJ6BMVNx3hdAG5
6RcgKQA4zDm9k3lvVRa3oL0epZQaCimn76QDDiT2vnHlK+6Y308JvNrP8t4D1Sym
xS8R8H1lRvKncqP6trjmY/vYt/IbcAbFOkJGbmIcCUIm+Ij2HRYIDI7sXFf3TEAF
QT93snCjIdZkrtdoJ4GsWUACiEF1vcOKXRjZEUHR/0pXjfrTYt/VCDlFxhtoghDY
`protect END_PROTECTED
