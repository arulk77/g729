`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAI9V22R0oxaXoN/JdDDZZ098SiGXFMim13uDyD4sqMk
STLkWDUJBApf39qJmeYXWnUWwZidtECoE+I3wP5Gho3+xrcEC4hB6kccWZrNlN0h
4WvBWezZYN2qm3NwuVvw1qTEED3lbswXuoVCrpryXlLVsXoPSAXz8nvoscSd5zvQ
`protect END_PROTECTED
