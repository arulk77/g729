`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xUW55Kq6kpfmwFfdzBGkhLvCkcltV2ZRPg1i79S8VY7
meuvbyBEYRh1od5q/xqp2JccFLOQEygwAndZCsNXiOLhKY7CJ9ICP+36Hqcs7iJC
OYpuccvx8FQ8jTjwJAk1ZaNeF+uAMNOCtUKejp401JPgua194HizWGDqtA5i0iE+
Zs8JutwQdFyUhyjhR0LZkbwfXC53nPWya/nvE35ayrYUmiRuH6AHeYIg8Bs+Xqpk
8v1OOVDtMUi9VqYjchaVLJcO64lpNANTENkqZwRrJIWpVypBUb16V7pnNgWyYN5q
vFvLRDNSQxsx+HL8ObliVbU0WuTsz1C7Ug3IG2mX+zNazDHhIdgJj1PMBmJpp4JI
ZOosuJtWX1y52fWieA++rQ==
`protect END_PROTECTED
