`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAnG+6+k2CGRhk+JQW8MRTxafeC7wK0EBakM5opGX5Z6
+y4/fGiq19DEXM+wqs+x6TwNwL/nImsuuqWfZJRD8QaN2KuURl2p+DI2+ri5msbv
m9vHnrK1cyaxyIwUpGC7p48bwJaF1UFP7UPza8zRmwAQ2oATcscNpP6sBAHWd3Cx
p3TBYxOeXuGFsyB80vLathZrX+aG7VjbLhGnAazst08huPIBn/LuNjflV84VfV+J
T06UEbbv7V/44dwmixqXTA==
`protect END_PROTECTED
