`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YJP+D9GYulpZjL1+uopbNJe7XnjzMZjtzk8JYspRZbdD9FCFBrwfYpbbleoHix7m
Vigs0WptrkkQ8PWx2P354jqyYY1b7gaXQRLISELoFdrGjCf2ZNgurYP+sdD2JHZF
2lB+/Nx+9DEagzFK7Fxut0VGb/6NmHDSHcvcWi6Ib8hIaY9bplp0RqV4qXpCLUd4
6voXRI5czM14p9IrqGKjJoTGnHTGY7EZNAzAQZpT6nTjMZtGyr2x8b6+XG7Fhao+
PQN4wwO3RcMBnYyvrJCtdD2uhUQh9QIYZzpmrTNBnQapr8fQeU/j200qIRqReKDx
IqNE3AlgqWxHifTDcVkEqG0bgjhntOQj2rZnmhBGtnE=
`protect END_PROTECTED
