`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCUTVIeEOQFoUlrmWuZU7cIVRGOX+3VECNX+d8nZ4tK8
Fs6rqbKRrFN8/vdlcqIxK1ZqBjzgIxELeHnEuk1OyOU/bFwvl2YvAa7ZQCqYE+nV
rjR2ZM/ni6V5cciuJS/B98954VM+GtwHtcrlveBNPp0svneQjaNcjzzopJGqc5rc
`protect END_PROTECTED
