`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOPT1Ajyq2IEZhM+3C29hvAZi1X/of/i+riD18K7dfYV
71kBc17PeUq6JEXbXZi7ZMNkx9FSOTrvsXlXJoGmJz5PtzpjY+wmdJno6YHZJ2AL
xhrhJdSoJw8Hm/aDMUSiLmvX8B87LqzgGXeqUHFOKY/ZA9nmeSmedfhwqE+5b9ne
/oCRcUfKOIzbeAeh4kNRSN52vWcDgvrxf3B8i431eJiXC6jQXEJmqjbDrUhtX7Vn
`protect END_PROTECTED
