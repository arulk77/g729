`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePG1gU/I2K/3EvEBP3oARJQTL075ZE7Qk6eWfYApkB+K
NPLCvi0eJgn2yqJr2Tb9Pv6CBwu247OMs0tpTjLezm4cdVpR1bt/oHz2mokZcFrZ
YJJLUGy0wcwqAYDmBqpE2QFfRYB6FQiS98dTbgXfWDCN3JQM+7MwXKpQ4zYFYN5M
fnjb4UCrPX6yg+ld68xxiMUhNHdBf1rt2wTruCqlYqDEm+bdHVLZEHP61BVfl8pL
`protect END_PROTECTED
