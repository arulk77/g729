`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGKDuxvw1NxuHAZfvg9qlgMMTx4xuHHUUSAcCWehufpW
U+7CzRN2O6irrC5P0T/r0yYb3knIXdrpMlvYk9NCa9TE+thPafEWFch2d6LzcDkd
gUmpV4hduzY/xst0hEpDNH3ZFy2jGvtRoD4GCVcYH+bJdg+uJ+ndHOLiy8txWxb9
B1PvjneARxHtiV7bwPBqkFT23Gik+R0CgAo59Yv6S+fNfb0JQv3veXwMuS21eJvg
0ne10DvUm16xVTpQFRAqUDAKDsXJW5lFBvu7uU3vYa3R6Xwg71HvQ5BJUIBnsnCL
fc8nCCf6FSsIkJdCzfyZY9ASwNgcTdRKk+ei3zP8U4KLhyhl0jZRnHrIVOxxqU5y
ggMnejvJknfwc5FSP0/ovDKKCBxOiDQIxu1TauZtWnYfzaJA7hXYg7zjEvGbQH+S
jGmvtCxdM14rr19fXYkXixpw1hdC3N++qXIRztFeyRO+KVGV/hpVPiM9Z/O9SlQx
obTgb6CaEzmRiuJ9EEDwO1fuWqqe57n49hQ+lfWGSulaV2V5VPAjKX6AVET4gokZ
VJaIt84pOK9yOr0Kevark+2qPnsOLB7oM9wRBizCvDSCqOhhyjcT2v60I+mz/69L
dMZwwmsKzowFkgeV2ANaGkhtfTKmpwgQiiIZdq6/NiuqYfSVE9Yn+qZZlqbGxBR6
UkAZTVtm6psYtLR7ZPKcsspcn4S6FZCk5X5YcArGFSnQT8u/SD91SvTGk9emeNIl
SVeBFcZmXjaqcfNa2ESqPvy/wyrMl9i5Qn0EJGmHQncEAGgYrlyywD77w2bDyO4k
gM79W4a1EtQ8Dw4DhWkYU78nIWLdMSFk5H8jQQfzmBAi/Ti7lNN9YUH5dG5zo3ob
M8yqrUGhGqjmAOvTvq1VhWPFXkeCWiKV4rIcfiFvoe1YLmPX1uE/jjPC6BMjWGCi
26866cDGERtwjdNY8urWk6GoxesN9E0xfaPO8GCv2FsRCVytrAp+RkP0HjeeNdWI
aBLXvqKGF7+BpRhVHgmT2sMXju6G2AxFsSzUEmqN9IjN+tyQcbhqfCbRvc5+6sTo
OSYM2fofsZrfKpKTwzbxsHfz5kNRjnuDDiUDiTU8iixiQAQI9jRZiJT7ejKMAFMb
muUQbLavX/1udErBrej4OHFfdgyTvAD/yv0SlXr/duFNThiyD2uJmhYn+WUbgdeR
Y+loSmN7YOU1TTTPTS5NupxwxMssXMaXkqAim6NqKmuRr6ynU+SgnQwBb9qHzdcZ
+mTlBHmkis2b86xVycFfel+RZOn24pqjXZmCsS4XOkguWqUrXlb2cPEyjGVTQt7h
ywzXnOxbUBkuahdZ4C6FoTSSzkVwizrhxW4rFBwFZnqkn5yhOEpFBGqcCIeOESKO
Sy10qd8YikwjrC0leQ97IrHe/3TljLUSnHrg1nxbJ4J3WmNDxH3RRH4PdbGgwpQn
CN96Cebx+0IhVKAv+goE79WV23G5iIzBjtl0ZIF5UjmG/05+4AD0q9/4LTOt65TX
iXkF8aqnw9SRUlfTQAwNbhIYcZ5imRIjJy1TujujuRQr4ws8ixLlOvkTU29o6Vip
rZYPZQZ67y3sGHev+KDPz3xXUI2fCYB2f8SXwtBBIox19k/xHAOXq5XweOe+79my
E5O05UpuFRPIUYsP9sD9GsZFmTTahwFJa0b83goRxm6Gh6yINi3KstUBrme1my4h
o4QiEy8vlRNX2271W9J/rxNXpp639bf14vdl0ctXaWb3fm70Q6sgVnUDIIOU6xrD
jR6rl5s9L//2QPMCzADYw3KdkWEgn4oY7ARFJvObpbpKJ5/fOa2GWR6I8NFmlkUw
wvzdt7m31RCAMmxjPRyhWWllcfeD9JS8o5ECyi72BpKhKp4WHY2T2lca9dpxrjAQ
GZ795hwy/x7jN5DA1x6yZPOdOyex6LsU8YE5HwOKEptGQL8wTSYR8kKrUhE3pzUF
hiEpw/SSCKyWeMuStlINwuRia2olMTxw070s9XetFy8YIy4UKMl2xgNDQiD1Gepx
abZXTkANbdQ33BexwPib88vnebiJnFz9/C8mpFSmQb2smpUSAt7m3p4NIqMU9SoQ
ZjHt5YPv4jdPy5BTq3AZ8JrbVxHMxhQXEaVC08fbjUQn2l+xdxAj/5xV5nX8CCrz
pW9o3zkX6oUBkf7aUMzH35nmPhyqDVn3M/k+pt3VtxAA+g1xBHCwrMuzkaP9U2Kg
TiOy0FPb+SvtU0hfGLbq4M5sBByzZtCnrourYxthDr1jtZL8s6AfUn6VaS69E+tl
xCBLXKNe/1+7GcjO/STy7VihrQGDD79kM49PCguZ5TRnsKlPbwa7TtFlRCg2vSDf
slnWP+C56ONWDjRaQU6qKJEs2Al55RypqTDYjrAKQV6DmYib5mQ5rnv+Nd5OF95K
MFPArOgL9qnz9OUOKwwjnPYc2lcQ2pthMu1T5973/z/Pyuq3/F78T5kth/phCCFF
s8MtmVgY3YVKqNCGrBhEHH3x0LjL/Jdxa1y+T4Wbi9UbpvbPcBC5uxZA5mCgF2B0
R9JycXNmco1ocvsNveKZiAwVvqdHU3dX/Ex6tBXrj+guv470fdhxprso5qr6QN65
Shd2CBieyhN3oMUXNj5O8it7DHACucFLHRKPdTyNqPhSabOv+AVYj6unN5fTC8d/
bHMTOoz++PeDwtnmWzKVwir8FGZTVtLEnE28IpZBwJ4ArPhMHOhvMnOAmVVVTjh+
AN/df9AYxbYVoYcN6Iqi+gJ0VqRg3/TDUoluKRD0LFPU9pbZVdEqMtmnlFLm3wWJ
vjE8wLk56eZR5vwTG+4iqXjKYcncn69KEhB3keDT99spv4+mfcZ71Rt/cQBtRRr1
8YKdXmVru1FZGQETpE87AvZ0FG5vbt0UhMsnzN9Sy12V+KifUC+uHHiLUMtmydpA
7yp9W8sVBwYTpQETCfgD0KOsc2A4xjxstuc9m1Hu47g9ilolIKppTyDnRCXAezbM
fyHIdaqCZDTm0bfx8KfDXEpcFGeXvqzGTXt+SC6NJQxvWBGSZsIsTcs0YLa5MAcy
BkqNtLmhaUNNKy4GXAfr0g8204/PfV8Oqv2Zz3qWSZXsPoiVhOnNWZq+ZoITNuhE
9vBzyPTPkzrIMn24CnFt8y7O7PV7maRAukZ2SnT/O4YG6JtgyHDZ+bQynYZ6a7b6
QJD0TaS3vWT3hHXwUfGIU52p3Hp3mCQWH8vrqj1Lt7VYJpTg3n2cg2BsZL3sisXE
dqCtoBio15OhNNasgzgefGsJAVJVzN9UDGL4o8QifNazJcRx5MAVYRqXoq5WM7ug
7JMEOuvhexI3YtZ71Opd3fzG4HsUhS3pMS2mW4ZSoYz79TxWOaWD6QG6azwC6+Xb
QPC8+hcMXiCL1C6KoH1HfGQaIgekbEUCIA9SbBcosaksQYeBEQLj69OP8g4KB3qy
rzMV7nKDWWO3nCCOP3qqJjBDyu0oxyIVVmMOE5QCe81QzvR2xv8qtrQ7jBl7KT/E
2XY5UysYPCe7/7VbMP2I3G4J/rZxQaKcKs1dJmi6H2zGYNA3oibMph7jwoqmdakt
kNg+gCciZKobgjseCTEwQYBIsEyWgPha/BNgOlZYNrmhu79a8vDbQjMU4w05WqFz
dSAVtggg+1A5Au2ejOXWTXM8B/oAcyf+KCDRSyCBDZMxkV3ukfTljWzuarrN7kh0
IreDA5pp1BGYoEWyNN0XWXxQDxMfAo99CtHG1/DSNdzn2SbFDzTZt5UnfOUwTquy
GEW3njtF8RKs0a8c2Gp1bu7XYvsvj3bmu/NhInwjOiZv21CnI4KVDhuAaJWqitmC
31Q8SFLZE0oCLSZmXtEfKp8/chQtxLN4aB9dt/S+u57XTCxw2s0WNN37Uf2vIUs4
ivsYZUjaVRQdDuyFm9bsXZJObKl5LULJMi+xjAdeOzsKlgE1MQG+ZdogT58M1xOY
3dxngR0zA2ZYP0yWwy2nDAa5br4jw++KyE8jhVmjY9/swLHjbO8CQhIQCxaL7otC
OD/AWnbgNYVmbWARH2xf+NPh6XVWsw2pGy3WOAsieP9gE3fb84APzRcksNbuO6+K
yBCE2mO3knmBtNO3Ea6XMKkL3I10cF5keapleNmwWftTKizYRR66tbDxdca8S3kH
l2cbzEel6hIWKWL8VnfNZvbc2MKM1wVkyNl+3zUGoW3vA+2bbvBx5DivZZSLNRQ5
vRI4fG2zlbgRdxqfc/+iqh0YIfdxQrUw4CXDhE+2/CvVDRPh4AQPRUcMjauiT+gw
J/o3FHXyrhbTqruZEaIIAqSTiX5ic7xk8M051I0OKnsTrqVxEw+7E6zmraF7I2ek
lw/+YzcwcI8i47Rwzl4fDDLhXTVvjvsFJVObVppdWxe1FhJZ8npVNFWPBCnkoMXk
TaQxxAk19JnodLuwH6bTAmQP0sQ9Yk5+GLLe/sxcPYLr8IHXgB+iQFlKjoltX0+Z
TURwu0yHBFBrA+Dzq4JWcn+Kw0PmNOEW1ON6FQ2qN0wxX+K4SmNMKd1GvVMwI08l
eCv1IZ5DM02UYmhMBlBPBNJNWJK+uAuJcm9k38EgxN6qxvg896RoJCJQzbNiroL/
qi4etbiHK4z4wbcGDkI9wEQl6gQSsEqleQ6KZHfcJDuFFV2uEsarVlNiB7amuumj
aGPQO9UuovtOYKfw4RrvRaNUGgxEX98b8x3BcK5gbfR2j/eMpOhsFyot64cSXAcb
r1KEtpx8Tc/xZ+qUohOLvC2f043fQAFJoxVg1Yj/fZUg0/yM/EvOYL1Bf3cYnmRb
xwXPtQ+IDq8FZEFVW2WYfYbcZJQ0r2Z4ICAZeCnDPCnMTUoED60xW8QpuUUc5qrW
x6NlVRVNOvEKMmej9iy/Eq/Hr2H1ePrIh2dhxndk5rFRXvbboROfTM+hegFOJd6w
tvlXEOGrnr5BuYvM/9GmidlnMpRpzNskOI1ckTLA1u+K1KeXexNNPc+9PUMRBP2K
NgJTghIPQYcCyjLRxeX+AR4lgYCV1wxlqczXWIZgkByf+XtuTJuDapENQnaSJZf4
UQj92Prc8dv9uGXB+EyiX4kb6Uxjm318dFt2LEFCClf4aycmYCFqQZNLw0xgGGXH
rPT2IR45wRw3nQw9q05VvfgF2Y/v16w8PA/9K6sq0I0LwFa5LQy0cajM+NNgEtNo
8rPS6ynwHAy3g5w9rr9krHXK796y5kL2UkNrpkTQ/Hbvo5jLdJtrJi2rfMwrecnI
7NVYE5p1q30DzwUHxPp+wa0r2S1UxTL7fBE7z47+aB89EC4QjoLZDiVgSsitwe9K
5r25uybo8TqjcYHsBzGiQ60vAnycCpsxvYS/E1VG1mXGwGTc7nzcTbwSxxyd/IhP
eRYTIbZ7U6KulHz8vB9FkPDhtWV7rAEkZC3GGsmfXHHUIdGrEXEtq4UoukfODn0y
obeoEGyFIz3pBLB78r4Zb1Bakfz2CHbve6cxk52Nd4CF9eDPtK7uehCnZ6A1U9JA
3JjwquK8oOovoHq3LlHacHYL3pQpEiU/gF9oomVgwnhglonpYVkLCon9QI9sG9dr
adQA/eXWd++iRgmr5z8wI+s3jITgZB1/0KAg3R4UdzbaavNDtImp/WYPLzZOSvx4
UFKGS+uE0SEfv8AJPiGQc1/UiBAfQDcp7wQ9ShKRyTWqew24X5ZEkVa8IvumusKq
AmQEHXtfTSpyZ3GMDytZjjaBnihgLTmC6nurx7/MslqCV8dRdtQhJYY7H9ZyNH7z
5VZvyY/7LlZQDhiRnTrTXB2da7Vg9MlICYX7Y3AXvTQRCsEPSH8u99YeJwP7LHM6
bvbSIn7pczZLlCabOcBS38FnpQm7DvGUm3FZkiDxljDNxG8deHg5c6+t2z2ynPza
mn/QZVuSavvFu6gNv5pJ8V9j04biRyCpn3OLBGkKrkfrWVhgo+lz++xWvZ474vUc
5kvdoKF5ju+ymJNa9Jg/aBlwRGBH/eJPKPCppThY8LOgcDLgg4VGbgACoybyDrRW
3q1s5EMYCE8zBqxTM+LdJgaavpleQcGwIyXw9hXpnJvQXBmn1s0q+1KReUly34uT
hAQZXPNPuEG1YD83cvhCZnLQAE3H0n3w7N+JHAX0sB3NFoOqNTRyhYQVqwLTCrz1
PGg6uVSTKEp/SuvRF2PTA5UuNUxdFGQSEr9R1qyZmFs4CDaFnsNju0pj+MYdmukf
nxZTwVILByFfBGO/L55eya4VGSpJv0FhLGFhhK9+y6BrVZejQGyOrT/kd4B538+B
caXMfLyydx16lMAQ8TnJyoN3sNJAtYRy6rxEwm9N7sdTat+dMRfKDiuHmngouz7R
CSpeozbfWacxCypd+y9CtX7FPaTOp/OXVJNfoL5krmtGardXbJBeP2UDKx7Dczpf
wna3jrRJIxb2WlUKgdy87CGAwL2h02FMHtmhLjxvoovCUcdogB/T0033rK8CSEJm
CgO2qE6XgTk0APpXCLprH9hYCJX0pYPJ2kMkVybAPsgas8TCui2w6uCUzWamXpUk
kN9pYq5Z/HDuFoCGftOuNxb2lZXhQmTs50/StslPkBc2zv5iVJTyS5a5foWd7MP4
1vjzURBEOAPC+2z++9hVjE6U+f1DdyboWOSGJ7VNgZV4rPI/V0b00NJ8N7mxzlrV
Ej8teoZc2sDZsiF21iyQaw3hyUeWgdjTAWus0j8MCl+Bhn4J5vVSaXFc8jZJmq1q
3gxBzqJnlpnszL2O8IOBXAaGKy0U/Uf3gEPLhCHJvq+E4hHK9IhvuuGaHy569wbF
PNdVt6AVey2CeJWJ4sjJkEh6zMpZi5XDP5CanvlRr0l8WUDbWbN5zFvEe0M2rb/I
yeHzWqeUkTL52FpaDYkTyGQkjbY3hJy/XWVDBVxDh4VDddieDpPHSLiOEzymSZzt
SU5d9DN7qMY4kAQgDemF5WAsvvEWgGUtj531C+MWwWmJD31LXc8WRTVR1J+Pt9E0
KuN4P7PA5BNS0iXGLOlsHqh8t1obl+cEqlFGtbENVZK1TM0EoU4iXj39vVnBNoK7
SYK4ZnmG+iiHY48vO51iCSNF8aqCJcwQFPsZBDwV5EWaH4dwoCcKXYPBDtvZ924r
XIzo2XWPeRWh7NRdC6f94l3ql8e9iv6pTYdBwp+4UxhOrUtlwa14wO+O8k9Bj238
YtCTagAJqwTxzy++FdLWklb5RsqbC2YO3T9zRdN32XbJmQ2pqdMiw3O9dCTwkEKm
Aix9ttFr6jpRYQABp1F1pN+HOsPyI7QMKMs/p7kqUmkUS4dBlx02abYWNiS3XNXF
X9NSJFagktSxQcKhrS+yDbO8f52vJ9ftZrXJRSIEK7mogzp/XjuD7IFHMr1aEhs9
KqZCwf/JabtznsZf/cdW79ygQWRCJlQBJ73QRREHE4UsYr0IGEc7zXNhQ0RRXQU7
0SfvhbEM723eC0YR0MIctF2IeSRVuVDAoyPSdAnnu8kD+E6Bar2gWZDQljwxa0HH
OBXQGWv9JDaThF+lEU/eOciAuP4RMfmFT3O13QCBWjamTRSDqbg7/dICWKQRnrJr
3FjRzO4zVU7TWzEKq2PDV+Fnnt3lnqIGpLg2ZfaHR/WK+gfiEScTPpQs3ZdKrNlS
xjZsVDnmbCIxITgr7NSdI2mwG8p985WxEeqJSuCYlbf9wmVULIYYNCBpAWUIFLza
4uVRcbMuwmqu8zpQLz+8K/cyiLzV7Zl0q2jkBeTXnvmw6r3etJoRjV9ZmD+TuwhM
JkIj//UUKJeC81JD0d2PfODlEu+Eb66BwOx8EZHzGE8ZGU1j+yYb2umRSVN/jfb/
dFpCZTdZcKblNomfALJnyYafjgdwGkn+wtJXlA2p6Fvg/5amvtSNwW4RXSSCyohE
LLuPN3xvlB1cuqyKpRXHuiTaZZD40/SmwYuzfh7zvgcJvFg2F9GB/ec6Zep2YC0B
S9TdJWcdvE0/BdQJKclNQvFlC+5NJFcGxxZSU3k6mdMjWDO7N2B35+ErqzOlfXxM
wb3JhpXmN8GswNWxTyiCLeF9OW2InMQ7Sc0lK3PI6iJ060ep+HbNbyxRG1K0FxFf
0t2l6pozZ5gef+opn4I0MN5kr5Xno5tdrtf0R/UhN6ZvZx/i4hAn5r0071Krblf0
iqMeJeWdtZR6ORSVgJlMz63OhjVJNFLCc9evInvMXoPihgL2s9HNzJdmDSwZFhoE
EFoarvoif3TlPooGoQQaBGdniZEhZLslh0jrnN+KaRBW07INb0+BXS/LfLZCXg+d
5IG53iVI8t8fRxifN4UZMXrG55V2FkgOBvgFCyeP9l27eZqws2ftovn/SoLwE2LL
Ll9qcpmZhJItX/QYUiJk1p6ngMFwDh03zNs9GYb/JvQq5aWqutEU3LIZGFbrbgzC
t5lLWpA3Rv1FSbCG0onNORrD0pPB3VI9ew0/Jq3srhJniQ7iOqGRvNZE/3pkcsz5
P0LZNcxU2O7QuqpklAZyVC0H7trf4mTcjV7ZJmYA6J4+SyaYxD94uuN7302654ER
Cyfa8F955ymke1UpPfGPEkfpNzjH5+r3gdbjNLYqeBe/PLO0aTXxZ4z1uqOjgWXy
bKI/mmQlhEZQV/ocV1/4q2MjtQsLz2eCo5Y2iobDDYdqdIH1N0YCT1Nv3GLDSsu4
OE57JfgMo7hwW/MtdaIMt/SDr2ShlessoOtroFN6mkRj22IDIWO4EQ4cB+yKRKwb
5ON09cy79gOFfo5g8qHxRGnWHynknkQFPQ2YEA2BquXqGQbhL8ZgxFHTno3vnX+S
AUpwuRH0Jkragq36rNcM8Xs86v/1LQqRFNcbsKAO6mMdLo0sxHO0gQ2lp0oF04Q6
f4GMiABc5hB+AgHtjj6l08jSbpbfjXXC1z7B9usjeudjmbNuP1oglC6uKbg8B0PI
B7dQb8FQlVAiQFo8/WkczLefbAHnnRvGfCdNp1BhR2gXat0QCKkLmsT5elGPtT3E
t8MkcQyX2zJDOq6Vh7PWAwiTTqEUA2k2OgDRfU7YaMbWGuPvQ8O3UUNkUBbezK5R
ze7xW9qaIXtY6j/sjnD0x1ZrqERqxEG85hVE7DTzJ+JFr0gxGUaDcCQd+z8BJ9uz
2WJV0ov4ND4ctuvARqScS09KQQXm17iIrq2B9NToFF+myLEZR+WRhrWAZP3I4PIr
ja63o0lSSP30CEfEhD3R7Gqu79L4dIfcMsEy6yu9Crn/m7bCrpysZwhZO9w15ED7
QvIn8CS4wsgxR3SdvuFnB9wTR8l5bpe72dNlZNDSkEZe9qxtyGxtwIh8iY1OcPhB
K6UsivWe0cI4j8lWuk/G77yGzdkQKCBd5wkdjYV0Z4q13WxLY8Il8ngQ4eeSQAd1
buz2eG3ixa7A794oicRFsaNy49ZRddeWSRciL+TlekXoijDPU6OjRpKKRg/gX1Fh
SZlCgWNwD7xZSN/AgWw9vhhhBwHHjE5uJ4GHC+Rzl4usJl8h47uteKxU44XyR5hP
xoZoLR1F/8CyeKB+cAVVoF8J56042hiCSMdknEBDCHi5XzfuValhXyRzsQKElQAl
uNMu6+a7jPYQYOPWRBKILvcJx3KgR9qquCpXmf/DYRHkckgAiLhzyYGXMHPnv+sJ
rr6ccKtkK38iWr/jWSpVETF/n0n6BXVEwzNKVUh8s27SWp3F8tx5Us1mo2UsQiU8
78RNXqf4RD5iDEcOfrtfVfZm3WzZ/HpmQL6eDDU0cvH5aZ2so73dvWOq7fxel50L
Ew/I9z8642IY5ow5eQnXwOzKmUalBNvoOjT6Il8acHsIIVoyIuvpuNDwDbL3iAda
2La3o10Q+iUvVF0a8QJ2P4yP9+PpclKhG/axlN+sVYUO7qf35pfsvVPE0eG1UHnM
zQidsFX8fKygO/0nu8V5UxfUY4UzgmGPpSXtrpToDu02pmXL1oPhgzFGWf0guYtT
nosOrJn4vUphnoavulYhpcRlPOC2d9+DDypfo7qmQh1w4wkFgewY/5zmje+VKVKG
wMYbAZoJXqy8tn3cSNch1PApBv2BJmu/1hlNrqaJVmzWsyv5mwOxRYPe5NiudUaK
Onc5PxR2Z3mVPcVoPIb+2V73ZXq/haDWcp970KwXTjJ+gTt5eirXteBNIdGCgjnl
rhnbyx8Vp0xRg0fYFMQ9/vvaIVYuxkgcykZoujhPrVw0u2LegOjfE76HxkoiZb5m
071eTkmYYSz372uTSmrFYxM4zX0aXELGG3/rHD8B2D6I1CGiqApUkzAlalJ4EcWY
ei1uTOnxiTpBGlkdaPqQGhkJCvhlrsik4WnTkhdLT62UwINDpUWl2Ga3T38oi8tX
ries0L+Q41vB68b3AXqf1DSRIpnQ8+xmTM3STHo8yKfkwCsgC6oVATFTdbEWQjlo
Gwl8gE+tQKsJMVN45FTKFFuqiln745BAwnKSb8/ShVOCTtHTCiVOdvbZq3JvsVDk
XAomdsbKylLu3ykz5FmDjENBt4/AvbE2V2WI+mFFU5yx7LnjR3MrQCA7G1p5VxQY
qw0io4rlvbuxYvtzCzbeT630YQhKhhuNcTU0jiSc/u/PfdnAPe2IUIsggoEzoouo
pchXY1F/GG3vf8i7OwaRilcfvPhtux4dSIz0TSC1FdzuFy7JY4nURpcmKfDLe8Kj
iNV4kOcIuqwmGokXRyBtPGfJnFrVQpkxBAtZaSH1Wu65SoKxhJ7ykrDrGruFl2Jd
g/S7GwOewD67RatotWY0E29CB9CzEJeR1I1PZ3E0j/DBSXc7EzVqPuR2/eD5vINP
MWPaC7oYx7ZNjNmaSaialFpMYH8BGJuQkYMUTvFMZNDSDPVIrl5woXhLNkspqJRl
Tplpwyuj+l1DeVRwg0d+yZ2+UKcRYn7ZPdgjG5H7M6lweoljqIixMpozWPNqGNQd
KrmOPgbCooBhKNC5EmSk4EfU9NEMOgWDX3t5vAT0Ab69R7JSifYDzzX9SQm1/oyd
e5/cBGNiqDy/dF48TzkAVqpVhDvrU9DUgCegWI2l8hOky6df44C47eGsvJBDAPtU
aHhqmfW3vhPkEShd58nlAnC+ohZcZ7jUwu40jH89iG8YriieWGJv+A5GkEFjnGsz
PbyzbeJoyp1NAc050fTmCOSoscicssMJOB5E2e421ji2YfV5apa+flXh6YH6ftCx
uNXz6OnsREmmos+V6GNCsOpMZoC/c3dpRn8M1C/Q2jJsx2iAQFVlO4mzEdMBeRa8
2zbNyMVgmp0i5NnAcqg/K4m8CRug0DaI9od3qgVTgN9isVtbokcUA/H/0Dfb2o8m
82tVDvE6fXJir33OgrAcRRVONezrPVfdslBYgkFeqFtvnOzo5cmo3WGILXs+QPO3
Q951Lv5fb98aZwVAt21HnPTyDOE8q4dqTBtnMEYMjscluzyJk1lrN0TAxEF+5Kmj
I3g/Nxt8Lc4MqfBIJFdHxYpmmQiKRmDmlX+Jk4W70Q7E9vDes3Itk8Cq0aDfw/Ud
itypPg9S8rumajICCGR56g/oH46qd1pwuaQrnUaa46N7NAYQmW8YVqp5eXVz+dW3
Zp0uTigbgpBQhkOusUaU8YPFK99S54EXT1DcbcAlM2L1xH2glww+DNXZaRVmkm9G
y4zVVSz4PY8CPXRkr3QcQB7Me3wXch6NlEmiV6WjLVBpNFYSipo0/65nqeWdHg/R
qRdOnkZsgI3Q5EYIOBIeo0Bq6MJspexoEf2lLic0VLX7xTSEUA68zqPhdgUbQqxg
8VbQT53djv50CclhneAXuAwKfd7d0nb+nSW29USIlTyXRg3E8KipJqiLKfU8mGob
CTuezqYPn6kL40mWJ5xi7rTXGnN8ovQbthWbcMN4HzHo082p7IVT71NGm+natHSO
3lwav1VRhuASfgXBeQJpjsdLCuJ4pLWhEG+WKMRue6uogi2M1xQ8U41vFGFYmDvx
u8X0fLhcHinSwHC4mk3sr+UmAwqVwj54KEzyRJHSC7LJ3tXlTzJG0+Dc6AFcPufA
FyjwinNk6kaqDBvkFLSaHqO0B29fAexgt3s6FrLhZknxXvozOZMj9LjbIGFsII3Y
xljd9xh1S/GNCUquzCh/a44ESBkg4fS6lqSByY9z4zxSAQLvRFE6rqVd/TuAMzSc
ToHI5+ZmZLjUmufi0tt1CvKngAV38B6sVvld2XzXXDxB8uPVii5EtgHJmhh6Pu/x
1g8N/XDqv9JU5kdjPv69+SzGCG6l6G0VpQBx24ajCsAZlLSeyZpPpcOQJDLpp37u
1FzOp/MjOet/l07VwpscAkGLkTFl9pLlwS/6Xyq16t5rTawwjhVXo8roRfkjzCXi
PTwUd3GbEcxZrxp5UU48hvmW9Z1ve591GPUXAlA8ZcUhHwjuteVdYLFfPzT2kIGp
e/2xmvAh0+bMum7Qz9OBRmWQ3iH5syrK4GStcKDuTMC7hiEZVLro/OqzGTnOWvSV
gGb2UVJXfS9ZFL4FNQXFhOgiKfwhafiR/WNrObEC/wpuFXmg2S4Wg9TNv3hB26Cs
/DZUkCB+E1jglLCp7yTpfcDIPTIVhFUZtGzZpu+nDDR87upJ3Gbd6SGeXIf1ZXTz
AM4EkMa1Z+WUfqkUuh3fPiLOIEKIJ8pTpZAmdOtud8Te5Vi61UKrvJjzrxE45fCW
pEzYMA8Z+UbSmjN/SrJ5e3BqHEyPErpmDnse7prpyoiAB7NeA94it9J5nmI9NZ/K
Nc/N97+vWkWE/I9wLc4Iqs3+DOeL5ZfaiyUN0q4DHanSUIMr39ujZBCpLinmqHHI
/OD3EN4t6T4EltIvkUhXPehWwKT2W8eb5lQk19O+d3j14hrnxyqNV6o8R5Lemh5X
byjkkh8IzkDbNHzt8um3oRpjKxtasckV2j7H//KhvliMCfo0rcboWNx/H3G6Hj5S
dT3UyyoHvzmiO0IShsBYC3RIKHlPiewEC7Jc9C1+m9xm0He2ovfHsVGBL87dtOF2
Ge1T7CvAZflVWKgZmys1T59I9/t+W5x1cYksefnP8hzZZ/GOP1TGa0pplanBB4OD
G1Yk68PjTKml2MKYHBtzl25da7IpT45eNkPzu/QguRMZBy83l/XWmRxIF5CURsEE
9F92iRhBtMqX5/++KAtuMw==
`protect END_PROTECTED
