`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44vUP8r1ZZRfSBEzGkSUYkedt+Ik6kvN/PgPOa8Nvgws
8Vm62HPAUjkPzwxuWeFo8LVnXkY5hmO4dtvBrvhc3mXMag46XKuwD2T3BWYHVAa8
Bmr66LZUNeMf+NfCPbY5y+kXGRaCstp7ATl/DmWTKbGe/iQshTJpxYzcVydY31RF
3RneB0JaIm1pI1v0IiePXLUeNYVXiaZcH041yH/s/Rh8sTCblhgeXFGp8eqskjy8
iKaR/PSaTfmcBKxSJf1v3cWnnk5q2YuRDiLBU1yyo+Kh8C9g492aome8zc91m+vR
llYU6OemBsHmY2YjU6mqjw==
`protect END_PROTECTED
