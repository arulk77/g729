`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOnTH8syDjoDxSIczosdOabfnXWnR2leZjteRd+eCqTR
0/qsDqkNUOT3A52JeNb9SMjYC1Ta45ubzWVKdT0k+NMixJh8EkphIqm6ba3Txm7t
v1GgSySa9QB4tZQCQxgzTQ/dEX9oNg7KLDAFeK3CaygLrtv4DgbokF1LwPvpyNT8
4EB33SULK/MET+r5qFjKPLlAgvuKS9igdPdG+KAYNaPA4WyOcUmz4QdY5tTlXlVQ
DPENLgHRmjvqsq0IQfSXsi6xocQbTO+hG/rlzY3bmqqwiAFWEdyOM46Mcs5FppUV
uHUJcY7vEtVkJHAC9faGwL5MUnprpgCB/O8rnXET/8L3wKrmCrRLjiG5s+l6MlSw
/0bHZlzoliR+ZNRJcSdCsUSnmVasBZzfwlO8qTc8hNg+8hJoVGzWC68PCSEnOS7v
nGB7AqF+KXZ9IZ0iL36S6EBS3KO5ilrxBKrGj9YMwm+bNZ1vwEbvBn6VQVNXAtC5
e5vc415uRIe3PqHlmHJ5EsgMfMu65qlwcrIFH8GgdiSTuFCZ+aVo8EznWQugye5h
`protect END_PROTECTED
