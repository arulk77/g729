`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CCaw7NjzpMO3fBiXfv8EvY3sz05AQOrZmB/9fzemgTfU4hMwladkmxSjCyCWkxaR
I9/fbqbpmuSU4E4vAspcvmaHdUqYh6ohw3NsBZS9ix5HT1QCirJDZverUwE/ysYg
EZOYj34ALmxjLMBpvXKBJKyeIrOiZGXPujYDyN3CbsbNplXgCLPgJV2biOQisWte
czt5PYlAh0wnV/U8fdfmROzhVfYaZVvQCCrFAcGCr6qZenz07IFiRh3xtOBs5JuW
Hb8jJE6Z7++rnPCAZpnntTLazRWtYpokqZI03SE5gR8=
`protect END_PROTECTED
