`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZY1vlwoEHR75Jn88WZwLOO5yFUa7qmCMg+MLh8CBiLb+u5KDBMH2bJ2zlOJGT+B4
I3nX53kn0R1GI8cjOtrsK7fe0+rsJ6cvPDSPxRfeTGaQRt8Z6EKHApS0A7rQLWEA
ZePnQuuo9fbxdl0QNZXhuEWVoK4taJjeoeFcQOw5mfqkh4gYP/vy5yvYKv6TJ82s
rwC/+XVtwL58F1QTnZePS4XNoYRPflUdl2RilkPOfkJI28iSgu4MNLW4S/ARLIEK
Sb38uT+cIGolPxUL5WMrnLnVkutqxFkXw9qFWyvw5nTd4ztFIfrgp19kNVJSEv7q
cS1jHSK2Sr9L8ynArqogk1W3s0qcGKDzqedPm7YsKgP+wPKUaqo0/AI5tPhr+o1L
SnGG2hlbDLRluIL3JMr7T8ZUVeLbSpFvJaduDab8sVe0HB8kj0snpOh2lYEX0iWF
lxONwFnQjTVhkb/E8wENZOQtgq3rHPr/w2RxmXrnqS5IMwei5SJmpyhyDXpta6lK
Gaws+hl1wnEkIBtydHvQ7g==
`protect END_PROTECTED
