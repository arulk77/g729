`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAUCNf+27hs6dh9ZZr/KNWwdw9/kbhLbz34x2SgPtTGAD
D4lsAwBrdoDJBFxfifFC1seiB4qikRDUXFj08avNUhPjLBQ2m/xZ38HzcsHxXiuo
xchHv0zFr8cDJfG7DgCu0+FtfaT3bWwrug0ucBWSMyMKkaylMhrFzaHV+dei9ZLx
kEv/gqESRmGh/d0o2laoXL0QJObmAHTeKYHm2f4p6PQebc0409HHETJ60yXAJP7n
TRALHd+NsqxsGwWSMs2VZjJFJIbhWBKhFat4J7Or9HWMHXGG7D5nMKHdhZdk0p2s
07Mf800z/XcLNdoj2GXOXbcX8ruelyvWU8nff0GaPUJSRLdCe/UOtg//R1RQ4j3y
z6e11rQjj7WZ2FAk35TirdjXrlquIqIdPGOtN7GkeHPcyNygQcvtpPwyqP1zyxm1
CbxzPCdS2+peO7uz1WVB2liKnJG/9IDjcOrF4mpWZC4GmUPariuuFzcm/lGJnmeH
kHQXOhgT/UyurZEs9Z0x5FCRfZa5gk0zLTFxchLUzfh4bL+giPYwkHCbXdzzxVom
gplp7kW7GFgoGX1qmCBlzkhf3bGWTVSdRdhf1MtNr2e+KyaP6WrtJ2V30da/IK9Q
/2bFXaCfStSVC6HewMeRm6eNrAAznhgeaqziAn39bfcEUJL5qCU5Vivf+rvOfOHM
MKgUK1e3y/OQ4LbeiBKsd/f6LABLyoEYYs6NYgWmToJNB1vtdQXCEWC1XeIEjYva
S5xF2lzl0eCNTkNuP0HVypeD9DghAI+VffFuoXLi6vx/j7vTtlsFFsc3AlUVw1kJ
ILBPViRP7VNQH7ojtJoqGD6eQPDZRYIL80ajTwOLK+hD6YQXobYfx28AmZptbAXQ
sqc33q1ikYuoSWrypFSuAqzHo6AM8PI7cGQfM7mnCNKej05eg5uV+LIm9yay8sK9
guE6KCS1vYnHtWJ1MAbgNHUZL3As9u4QuvMgivEdi1socqNOkiAVXIgVKgcoQdJ5
eikZYnch1eB3gg602btfm/sh0tobHofthEYPm18lEtZ2JbgkvEqCOwe/5xqwkqtJ
0PNUSR5n8tr3I1jKwbxPFPSjFK5gt055mH8jsRcM5pbcvNZqjKXFIbxjNi7G4eEN
xs7WOztYI943SqAi7iwbzoTusXQ9zZEX3yxfCZnVF+uX1Vip0bfUecLDGhs3hkxF
o4MNkJKX0dJcN1jRPPy/+/A5xcJztVGcEVgNZ5dlBc9CHR0fiMUlK9L0Bm8qeTkN
ziGNgwK2J+SajaJbtkfTMW2NRYzl/SNZX70ysD4os4hsxrI/SkCdXPgnlWz+OQ1o
4pHmA2hj4yKwbcQzuATmcmtoJ5dVvoB30eIupKybGxRArWBg29zjbt8bzHBDDMF6
q4a/vLss+aFTlFFRHXj5aCUmTmRNA/ecI8+oo9y3C3g=
`protect END_PROTECTED
