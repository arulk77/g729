`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNjkwgDwDGi70gPvt5bs6ajcZwQJnUf/oc58QbEiK6zk
KvbvFeIKpItwxlwO1NYWVHzT+qkaCP9z79sM5wmEH7ntG4ej9N4hpLQZZpHqPwkD
JBclbGlCGa04+hY0398RdMYu+2mKhkvl811Iso3GgFlAgblcPMhKk2TGmqJsfijr
mxF43Zp8T8dAGgTQ+a7Z0bxhnjwH5e/BFfDEM1qbTO3iArSPlZrHAPI27iTGEQkx
LkrH0fNfy7sihyUj8FhHqENKjv5jD+Jzu/6eN617EazzmF6MiIYWyAdkO3hTz2+Z
qMq2FKGyxKn+vqvqll/fTmnjkUDriq0aITaEihWkmmgsDk+BgmoLYmpy6jFf3CbU
jxbI/vnXlCPE/r9bzb1Eb0rhA3KP9iMV62jyrk8y7e0pW5szeD/V/b8QGbp2OpdS
shAVzcazwbtwHru1WmZx/XeGsBKWBUHDvZzDqeN5WKYATDjXKEXFnHxL5ASXC/pP
Cv5NuI8UpyZf2J25kyK+4Lhrt0++oNWAcZH6Alc5NuArMagC8GpmQa/M/7Q/a2ji
Ue3B3dm+3CJ5JkdlyApEsyfELv5rL/+geMe4G4tbdrPxxacid+eBPTy97aP5KBCJ
oAseHKrsC4aoFUxb3P5qrUIv0sL08xFlVoS59Y1WLsfxeaVNLUtmrmprIhW1Nwrx
/Fps+xybQFO4ej8+519zP3K3fplBUxYzcLfe4g/UXDJPC0RPiyi/RQlkQBJml8/n
LGf8hhDO8tg+WoLq1AEkjDDTUxgKqwhwDN6I3rEPoZaz8y0Hlmh4LT5fiw3pCwIa
/G0/qRwmGzY5ETwpJ/lU1jixoblZbk374Eew0HZIRQWiwjwvYMAGNNnKpGBAVvV7
yXMG4b1UBuVEXoeQNKipcK2GIhSJWK9PC6G/+Ud2INlQupJo0yf7QUDEKTT+/yO2
vSI+jlTQl9U9jQa99vD/wZlgC9abEamthojIFouGYfbM1BPjs+5QjPts977KTYvB
lF5XQTKj4NeSBmmmopLqhUYQm46l5+hIRcyYy2pN4wmPLuiG76JWMFX5oKysYNGW
/CZCnBQzUTjyOOHuL5UC/izfqTZ83aJzx8R5cCkrD4ZSz5M8kmchhSZzGc27SqT2
BWrRkTHPl9RO73knMD4xkQ86oYRlLB1fWAuQc8kH0SR4jFa3Yr7gCRU2PfwCP61m
II9PpncD/Cg/fTKswVajb3WdQrwtCR2eAn0ZN3srjmFLHLJ5RK8bkp/vLixGtgtd
jmDE/7mesfYm/JYiR9dmUgOo2NMI58BuScor4WrLf1ohgTEb6jr9E+jKG5H1ybgV
ARYGELU60K1S7ISvnlYA7oh+O5RoPxsvES1RiVZy2n4O+MnWdegq5mgLIoCnuZyL
RUBh99/z0WwFud/WirGhm0U2bMhp7m4JRScQT6RyxFyui7dQ4fLjgfAB9cM52rpE
L1L899iQCK14FGhhxm7fV2n6Fh9y9+0KXggL3mArvJbcOxSfX/Ls+5OHtV7RW+/V
a6WTtXXdg4j4eHQdMAUzjQE/RWfTfUdU6Pxcl0iJQJpNQvr8cczXTBUlgRk10+hq
4BFAZlPu8oNPxj0f/MnZhzjGShLw6s+8/B3EXPyGm6g2fMCavqK9jW0RWUOKqlxI
qew6kB0a+DUrWqtaXFBgViAJl7LCbnEP94s5CEntG9krjUxYgH6eK7i9SAT+T1J5
iwdq2Vc7fy3OsHyNAdtZTIDJof4nykGwmJ5zzUOdH1hSducyaE5FkA9T0QdEaqT+
r5W2ruwgLbH3jUrL0LpNvgz3/u5rLu7GO/P5jQOSbB4+hziihpERtVb0htX+ILPk
PMwamMvvBxjuvU08ZjW9zEaEJRNqVv5kV18ipjqeULYTuY7ldkz+PBTE4+vCeZfW
Uc4aImi+VoLKtbBTJU/PoW/wa2Z53Pd2UW40L2lKyCPO4Y7GzKM1/Uh/jIAo+x0h
AIG5jx0bEWJjBMtVoI1dZv/JoBeLnUsXJTIRNjzyRN3uZtYpFjXCjgQKhbzCdUf6
pe2Kfzq5im0aLjnCJ26kd33aTyKLDgCsofXjniRotl8ZCtutsSJa3+2fU+o++fLp
DYPDt0sndrjhHdLd4TOfuH5kVvM0ccvzg+cJh0hpu5A9bj/6FpWnnjvoZmFnrsL7
2evxXqqb+diXVZIm/S+gFUr55gqMqxQUrcUotfgJJBKqI21FDSq48bQvCXI58ku2
LrlkWyuoARLZYIkuWTxNtscKcg7cZF5Bv+7fpKRMDPzm5EZazI2jUlLCXhnN63Qb
YTq/HuSqblT7Mz0ATDE7FnqQKsxuHfQwCKnMI0dbfapocBwGVmGIMsjXp6RDYYqt
TGhCV6d88OEl+GFJwTN15ZHdEm/U52t5o4pHr36iwPUWIGUBgGjMBdd8fNSPautp
/f5naxvMEIvo3tDZhts9Wc8WOdpiXCvyzgYpVRb2+/z2bgo78qVHZSOni+m4Oq6G
bf44BOlE302XkAIbCVpZRGx0otSbevVXQX/KA38Fp7gC7YUs6LKSFoo5o6BG/PRD
7nndVEA7hJURLy6BLJvikSax2b6FAOYw+iDmGOnhhNmQ7bZKLn+nBVndhds6sKTf
FU3y2Uy+YGw8fgVWh2pVBgAcyWlo59IxRFANU5RNL7RFbkivSDd5j/hD4/NU2Z0w
u3KJdiriIJzSC6olMJBptFNhsDz0yixyd0ceSxvWNzWxAJ59rAq6fWNw2NzwSiDA
oFqn/vlsxwsFQBbd2bIrVAB6wyPmNaVU8TKZdF3xg3d8aCWqLKo53oiZqJK2G0xP
qABjoHJoge6e3yraIPCdjmQzHc8VaGjRQplt+Hd+KljNBvm9dhKjVPNZasXxUao9
Mgs9kV5vq+eDaxM/hoQf3uPU6bee2NEkf8EeP8kkq6vth1lYLbve5Wi1VeAn7ldn
Q+AcLizLxW25nA4ceiijaxCiTUBG72TqHQBeryZ8ubr0aXwcmKtGuM4nON/idGdC
x2OcwHWSJhg+a/kJhltoBSMGA9V3RCp0xw9nkHAzRv+glCNApU6v3kdk8Yn6jsKe
Gwbphnv+peW6N+WK7AXq/vGLBbKwNMEp3dyb/aZeLO797oZN4LcIScZCi+9BhHga
XDlSLK+wjyzsHtwAjmaZMGMQm7cwO3a9/FNpe+SruL8tBzEOsG/Ias3haoMUVJbb
rwnrKb8GeXX6XnjfSIAQM/hIuMdkf/q0uV52xV7SXmpOOZDAO+uqVPPJkQ7+jQpD
4CcBz57Yl9JcjxWyemStlx2f2l25ggT7kJ0KPN+TlcQiNhQNIKsSlx8iZFPsGrif
Uqpfsd6szSn4rPT4RKrDLRJZDtfCj8z31LnPW+dFFf7HzlnXsmOdKzt6uNT/ND+w
4AO4NYvvMZR0u9I8NZ/zkByBvUdlJwgeEHeFOepeWymtKyvFxWMNZxRVqba0z0ux
I/QX/+MzGbrYZD5YRPGqOgOos75nS8yPjdMkol6tW6eZStP9SsjMUgG70wJpAzhm
/++YXV1+krabgXLMftayX7BbdOp8LVHOlXy12gPUAqHAuBc/91TokdEuW5jmVO0m
/JXNrfZfH56seJiCmQ1+hu77hleXuMdr33VzfsbwqDJfEuhh66z1qRVksvri7+Db
9JtjQWrQ5B4VLvaB5Ea93Sz8Hlo7PclN3sGnsBtx0e8Y4VcCaJSwizvMiJzTFCm6
RwKmQdhCKDggDetmR7JXAcdeJMUWSa30WUplyibUwtZ4wXQ7tb9LL1ib1dTXxLnn
86v0AuUsT0/95FdmhgG8pN7NOhhUD3b9WzJ8DWYQ+BuDcMFlAZTK5zhLJc5ELaKt
rQgaLSCqbB2wg4wxmXOQkgAws9BXv72uwid6EbBqXy+IhOXRw3jxdQ5EDh8Iycdw
+eLzU1tJRzO8Im1t3l8wKaMBO5pvO+hTno3M3t9u9ZC141zjvKeZiW/78tKvAoqc
NdS156JL4d8mvKu7OAn92mdUXk4DqeptPWfbFJm05Hdyl/zwyxWo5X1rXtAuaq7T
SGTfNXm1cCEFzv8Of/37kCEK/eeT3flxTqkWHVhH1IoPdqd6rdqtTLUeBOM7VYoC
ffUt/mszVCHLqQNzHETJFPz5IINFCi09croHM92zAaNJRJpeQ2hQ1ftD5yZhgwEX
i8a6HDlMv0GTKGRwBbAi5Z5FPymTyrmKNzJtfPFJGXso+z+XmAOLK2cIN9bNEyT4
SW5JygvbwW8pAe0Nq0t5Ag+wAMzm/tadCkASGigez+1PsiEBjvBrLb0Hjyo9zfuh
LfSqpyECHIJRWuTuCGXkgOzgTcSrOVLnSzbN2XnC7WoamDUoTbGh7eYOvd6ShXWc
qJvRgWo4ZAVr9atvMPq7d1IfiQbkmUpy7s/3SKRoTRl1cWImvFDXNqRwQe2smKUh
8KEWa3nopOgGet6YdURMYNyBDZQArN1Fs/r6FUWRS9HdAFIBI6DtERJQxSCCCHh3
Rdy8I68dMQFkgmBqv4kmmlAKcacyvYj/OrQ3MAwbZayyWuGUsGOE8tfnnyojgII0
fOMsS416tN4YUK0Y/qHmzuy7aKK1pz6c+AhM1UTgmkFZ61q1ZPiZ6LSxgLS+29va
GT+Va7MIyApx864dOOql72YLZfS54bXoKz+sL7gr3bukGXK000zP85IGYH2hcCul
eO6NnmOwrSJdq5ZmVJcggtmBdQ2CMCxkdOz4tP2Wfv0VRJ+2NugGTxp3PS1hy7wF
vrxFh6c273IQ7eK633ttcru/n9q+2QKa203SXdgXy9ahNFVP0FAShD1lV6KSbU93
9ErvI229e0GaTQQWVbooCJlHakyWTaJGVIMswgFByc9nfQpRci2ujwSEOZTL8qWy
TH+lgyBRTaMX34jx+7m6Dg==
`protect END_PROTECTED
