`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
r7s+uhjk+Yj8dlEWFCQto7jpEpzET+0o0HIigqRPpSYFrESJGrR27NbKqdg9SmqQ
HfqPpC0sbBMBwmjB8XBmZ3wKLAc31jYbjQf7AqZosUdtFNRMbQHjKrJnbx9LzqTf
GuNo6uTMkP8V9oDtwQwTIq6fQwPaWlYdSXIk4JUvQhczeOU9VMt8X1VZSLoykuFJ
g0o/CH8cBEyJDsDUV0OnPspmQ2PeDO47k1cuDmaZKmXmHViACVja7YtEpQIJvxJm
ErxlAUoPqpyPykxTadXQQjiZRAl39IxSeLfKW+1B1l6hJiY45+sF7dKImnxghWbd
an97OtaseHKW3EZt0UZuGRaH0V+0Bhf0zqQD2sT5rBquE3iboTJyQK+Z/qfIB8ZI
9T0a6F02JZYSAZSZo7hkcvlvuF6FQaR1NAI7cHmXKW07SUYxU+aMc7vss96+aUkg
I5LSFNYihfThhtEg7RRJFgitgGE6RziQBldixgtsA6aAGZ5O1/wVisB0iAySXGlR
Bk4X92qVci02dZlcAlrQ8+yjjYKwO6OkVkfhLEPFJcnk/gzvAE/l4RNZw7f8xDlw
s3oEAiw35PFbrxVU0oBNf5gHd12duPp/jvO7ejapsb9ZTqUzEvYLZmqZNtGX1PZd
c2qwGVSl+jLaLs5AOchZC72iphVqGA6h4rfTrjzP/zU3v6QpYEzhaSX4HRyi3crI
z93j4cyMgT9HRG68NfXNO55RM+RuIs17A6p3bqWjzFi2pHAfILVWV6MIhq8pzU72
kPaNnMXbWQW9fNDmTq2m1+4rDHJt4io37Pn7Ax5RqBFtlFIuM2kOruCQOr8TgyJa
uAcZr22UJxPaiUcEksZmS4yXx+X55bxYQzb54Z8xwlGjVRyHpdYemozVzH3gEwXH
hAXlciyjgysFv73WMLnM9kqZuvWwoh4Ar2eoZ4pJx15lF2HtLk4RT/R2g1Tw5rKf
5QDtmmT/Fhv72uazvcPddHHsgWsuMTTcSgl2RExoyu70O3JxCAYxAnwrSlVUjWBR
3r9xfgtxa6hRBngaoZV9huIb/fvlfZd0Mxr/VLleEvKYXwJa+wN06JhHYlbg1sGT
ubbGuzG7k/N4sbHGEIK2FD0MTTkMoXSs9oJCRBtDOR/gAzKmEMHIMSEHM5lwqCEa
`protect END_PROTECTED
