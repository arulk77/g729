`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAB7uOBTPxKUVeK3G5nQB3SHTmSEURKZ4TCWCyJju+ay
Q9HQotqbXB9CcRCKl6FgSQFphhZrjPkJbyrUV3QDeZWZFpefeZyObkuwlJqTd0go
hZKrP2N84KdWMkkZnL1Zf+Mhv6oQtO6QdeSYBLo0yeZvD6dZanV4u0YX9wJfolbl
/HgvzJo9+M5h0jT/vID1V8AMKL6pfqt/IE3k9TzWgpA6HRoC3OaBdvhOcju1KFZ+
AC6UZ/3qMfSGhocc/FS6rUEu4rquesYHuS0gH9AcRtbo034nEzc/0DSxq8p6ZtTm
jAC04XYG92OxaUwPWhEGUJrj18P+acN7P1u8EfDIDulmceYZzlB9KSbDxXnYWC/y
`protect END_PROTECTED
