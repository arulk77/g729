`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SSQn1QoD/Vq3H10us4nOPNurKSLeByR7p45RwJLfZ/lt
AhpjDpOjbhB32a6fxTVXogrRFG61DyKvX8Yf0ALYxi4gz8DjM8eo/8QiEJUFHSL+
NycMEKtzOfTqRpPQHYlYRop1/ibUeP95+PUaA4zrYfdTpBLGw0teKXafUwQzbS3O
wwQFV7LQ33JcyT2b8a6FxJxehgyBmZZIf3pPQeMO84HHuYRgZt9emGf28BjLZr3J
dZb3tHhX1tRpyR8E7pEBsWDdafc/1DJlkvcTgzVo0qg7Lzo2eVSeDAUqmhoTU8y7
qmu6nnzCCBs7z8eX5645KSUSQC3HkDqg5D94BxAdbWeFGRB2CRNPdEOtZOrels/S
hXugGAUQOEBGZ7WPLVYTIe9LYGeizgvtWHWuCOOQGvQQWD/43JCmGzl6l3O6LCol
VnqKN8HLbjYQEgsrxDnDxMZfWBv2x7dTWgoH/ZDIlOOxGdkEiImFNK7+rRw1HosP
KC6uH6a+NieSMakGceJMW3uWiXiIakLBnRqf2eI/IjOj5B72q3aq4W1acnhxXbXX
I2+u5O4RRp04DHiQC1CsD1MJdoxGSRgXXmqpb5Yvp4K3gsLlClL+yaFbshTvS0Ec
GdBih0RmMSwEdNXA/IScrZ20bYYM9KRisz7jrbf27V1VkulPAXooRmrCSeAw4IEW
6ZRLLiQRiy0qPCvkPI7dX5Z7fDvBVbGfk6nZIUNErsg9PElQNkF4aDdl7GaYeL4T
d8AcZPnGc1X4XfVUqT1H6v3rWb9LvHBWDzQ1kS+iqrPE/z4jZE9jLli7TjSIKf4R
wWURXuNQ/vmszNORzi3svAz6j2W6lTRJxvqS1hdkZI0=
`protect END_PROTECTED
