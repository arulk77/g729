`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBTq1TWDeMph2bfg1Zd08MxFJFyv26YwpjD5t4ZrZxrD
wUSytvQ6NAQ0GBo9QanPx4JaQQAkWCoii3fsuFL+rZx4YSvhSmnRuRF+jO8FL0J/
xSqxKqqyHQcI3UnESaygU/7i9dCbgMJ6s++8HtA4Dg+Uuc6axEnS7FBEtXSrprGW
j5//T7cQv2UFMbOh5X66TV24SxR26D4ztbu6if2swRQRpQxMZ9s70zyrCscmqLRg
vynuIh23mJZWA0MjNMfKtNKD324nHVBA3URm993PZF6t3fi3CEbd/rv63fmW7pnW
58I7crDnSHWVsksdjVIScNPdNZCWcNwweL5ofFe9spHF2GBFWZsaJLGKoL61Vyh4
23qVeE1UlAxcnFBjnrbHMobOy2fIcyt8n3ILfLJB8plIFdXoYlVYxtgKCFSq8pQA
k2WNuDBbFCzlziO+2CLYPrb5CMqbyuQkJwvcYhbRJ2OjO2AVWTjAljJ4aomL25UV
n/cxlgp+GWO4AvrDBKFuqdFz+38KwEJl8pyH1jb8Bz0XD8GN/4NidBF5RB+ThMD0
rvBnGMDGboPjCmGOv2Ed7Z2TuIhYQAtZ2jh5LkfTmupZy3L6z5wNJlGyRSm27/rX
PPfX3/vJMepFzGsH/RiNixzuhRZt5jgdlo7RLFbKs4snv4ZEKbXG8FNc80ip1LE9
p/O3LSiZEIXtPwrs5nu3TGtDfln3Ja0x6zMhsJvLHttPA3dx+jFA2P9z0l57rW8B
72ZW05lhO3N8UVAQaO/0gk3p9gWvJdW2/xnV2yLv9UU6Fdp5UYb92W9tpRddwIJ5
K9Km4rc3U0jGdzgdLx/a6cVE1TsxAYl1FVBE056IdyKibwYuLeiMW5qNOqMCPkZE
UakKBx3g99jrf1uvtS4jBzrloHof8fHOcUldGasYp9be00HMSfIeUCoOzk5qgoX0
KdU8haIb3o801QBwJxFLjDMEfhOec/DY8AQF283lfnYK0k/3dGM6rhS2RxSM5ceZ
YNLjd5HB7Rsb4Jdq7kJUN/pc3H64dojDjD4OovFxikmZmgkYWhAURKI8zIsDo7VG
iOCQ94vz0MDkvjk+RA1hY2SO6G7owWS13mK+n4TE3qk3KCt7sWFzww4DIpTf5drZ
5JHFscq3VxlPHDWMXiFZNeRCVE8Sahpdc6pQYh9hB23CC68eVcfeA/05X/wjVbAb
NWlM1czY1LiZe6TSRb9EXUmmHZq5heSbsPuubNALEq4yd2wZ5FCxR/LnvpFmzvC6
QkN++jqc7DAuyewAnZYdcsXNOaxnVNuewpwvx+JM+QkjHC4qOyFNiLz4Olotimyi
lE9S8xenCWRhG+/dQBqntzed/FGQtzanamagI81+MPRduzbGo5KDbuN4cDgAPsIF
iHuXnSk35+Cp5327v/Ez+DkrliI6i7yU/fJZlaBBovvE7h2D2s5vxrwv2hG5GKvf
lNxWcorbzpW73Nf0sI1uLmTD1l3oknoBtP7w2y5u3KxoKFzumE49RMxxe/NjOBmE
gW8R+j9iQZbv26BL1oD/4R6mQ/dLjUIQE75egtIne1cN/X6lr7QyyWRzZgC52QC8
oZxWSzjmNUsWJFOTjXueoYEkOABRNKmSddSLnKCpPn8t1H6K0CGgLwuQbsBW6ptH
rrXudTDSw2cw0jhGFMROHyiVcsSPjFwZnmtqWhKRBTfl3DFM2CbRAF+iU8lo67YL
wLr39uH0aznUac2FrfrtrjNaC2ybWzliVFCn9lsBlO71cKzfTIOamQKMCaWzd2dB
yHXd53fbogiVQx9folyz9vVN+W06N+doZM5ArBuT6vLCxfCUJqBj0ny6Rg0wyots
T/n9+Tkf3bY1LjkxQl4pglQX9sR97wtuBKy6IkJDjyG7+u68gw4N2wug3oRLvL+s
e3b8HrqWYgpNhQBlieMTXD085yBvFdviQiJ/CLRdBiwcTtD+vGX2c3fFN7olZG5B
HkBhP16WIYCEb3hKG4QjZDXs6oPyxqB8Dwi4TJlL+ZiR8GDCyy445dWlHaopxI+E
FI7WSHPdtitZ/bZrtjR0DCKfRJsaEgRNkTw3izIkgJXLIcHp9s7aKWQaljyvvWtN
1JY4oteN7TJVkqiQ+mZbbfpThwdcdX2diTgJ9rAJovMQGxWKNrAl1N/899q6UvNa
bMdwDzIadafFbZoCwVwVMOO1OLv6AXSpBH97xQUGD1p9trHz6S0+mF7ZeYnYYaXy
Dmug3fVR0nK+HAU0Oxg+oN53L1fYhi+bZroxZ67YYUV6PnAgaP7cvLzwJDTLV/QN
+C/F76953BipvisLy1JjGC/AFg7XolIeOQaVQqivn5xJoq+pR+RJM68GuTBxQAVg
iFRfe9H31TGMwlPnuCb3MhfXNqoAzV3kl6smSNpGsUe0P2C7MtB8dCbJg+NSMJXx
fiJEf5h3nuJCfaB+PfGRIKYTpmved0GU7SWP36LDFeEcOxuahVYAlBI+GWYtWhjT
nC+py0wyNCSiqySEPL5SMC1cCI6E/2IRxaZQxtCgxvzvPA4XSK0hAP5/vHWqZ6rw
hlP74J/3S2M+16QFCe13EQdZ8/wm+3flPoeXN7gionk4gVQBFk9xB3gH/8Mmb+n4
2Q5C13svlPmcbRAU5fnKbO5opp5yYm/1d4EJOs6rshwK1u+WZJfHU2uZSE493ifn
BZIqcXCBkkyP/Ygca0lgiw+HFCFnoOLomvdLQxTDSsC3p4VK09crlQ+sGzqSv1nK
9WTXozcsTncH9AbpDVhMhKpw32prxYmwlpc6F0Hxu/aBpXqmj2yDN0mu2e0N72jC
2F0fKhz+QOuDZ6i1vhbcHFNDtC9xqyc8nVv4iakkZqZIWHyYuPlaSl2sio7IqJ8F
zDKtyzFire0573NIwNf4CvDNY/WK2ug6JzXEyiz0C1g39esDbAQzcal2NyrqOqde
e64c/TNyIfpg1fVAbGg2Tqz4oKlfFzFvzM1JgR8QixdqqCsgDzLC1XLLTfXc9djL
vhAdBNdGLUULDQGAr4+/u4ujaYaQdfzgBWueOV4Jgf7sy7EIktEfGbAzWyqDsD7J
xUaRV07vQgz4L/Yew1K5EQ3byip/BgCzcQY0nVnlVVCaX8arnz6j0MJaQ53P5Ze4
HdiOeoPx8L3LiDOV/VFUEYBC73/brT/8kBPE+UTysWM2uJGE5rLOeJEaI+ra8YHh
8KyQyfj+1dPLHyI7oBGWbsKZg7+3qVPFXkPIWUTe4I4vGdM9i9nYeL020gWEWxrX
Q8jtrG9xJ1zz+ZnpNnKclaHwCYd9Lhied9ovz0KFQPDJ7ozaXIa4IcPmyjavKmZ0
v4CPWraJ6gzhaIv9G+5DjoImy/h4+ZcTfhpKuf/GSTAGVQoes1utaNM4NBYI/yGq
eB24cHb+k1uAi/uOxeP990Ats0P6XK5T2A05ED5l/H8etJnFZbwaiP5MZ60tVak+
hrlxZtQn43xSW6+iCNP2ySO4Df6OjOFXOjhAlckWSKz2XJ6CsSM17iXBYnpTGHPI
7O1UWyTdg8tkBatJBVnOgDzFoS1BMsha5ogTaDtl2J5/ZvMU59S6WgXTgCArN54V
rHFmHtPwkiSa5wg9y1WbPKk2R8Ob6B0Ff6K59rQdH4azhn+f2jPvdKLA56OSnF/p
4Og1MZfH2Ss73cwGkfzSjrkjSePFtTiiQkVcx1IBB+QgQhsoSozgrbtD6+C5CzXQ
6dMcXVmUM4NlTCg2ZBiBrdrRyWkJqUk+tM8wyN3TVKfU4eQXL7MCDq1QMJ3RZI37
NZZfWqXv0MS8EILjdBYWXdOn9tAGS95X+mSBjTUob+Xfmc/Zab+U2GljbJJw2DJ3
jwABeAU0tE45DjN8xI8JxaHSiqLMebUz+W+68MiEb1dB6bG4c+aQW/WiCGb8fWYo
YKcAq9XWKDWoT5yRSS9+FB05Msrpkedzm3+p1BuMgw/iwYaKLbz0xDgQkFxtbxEu
bObaTbl2lsfcaALo1a/9Ozz3pqIQTYNhCoNQbRvnoSxgQYoNzWOXewz7tdTmG3u+
SmpR4XWk52fjuuDSFaDPQHYmRjdsqAorGZNMH4nmUCQe8zJlWtyFMdkar7RC3OOR
HbAAaO7HhMc+2oAHb7ZfXGeZCl0M/7kljGxpccuxBkjLkMT3BZXhAE/4hZz2wP52
Cwk6cP+ogEmZtZs4kSD8SURsIY/glRQtTYDSQZUVxjliNbuPjoMaIJkqjANDFbV8
9s/oEooT4aPuuvFUyrktXrtXgpauH6bDUpnHldrXj3RGOmfmIKu4DmdkAzh5lcV9
B7+XPNHiuEKwiWNwB7QaZ6FSOZ/3TB0zXjDrZyXtL3odJxthHpIswamxbQCMg2lx
uezKnEj7XJrUr/ptPOSVx/JvhAfjpb7awPb/eINa8gzvugY3mh3LzqI7GKwI39ss
bVFQ5WFs07+C+mOultgjgUypCFoOPauNK4XmwSuZC08X/CTji5rZCaLm8X9Oo8PC
uA9Ywh/iCrIfLT8+v6vT4YzqwE775ukfcSs7j5KMNDrCnsj7YadUj94Zq/w1SE52
w5ndNtWokrDmF6iLJcaTOx0ygxtpZ7lJCa7pTu7j/Pb7qlV1O3267MCc3ReyzSBg
HZyZ25oV8qcEh1ld+s+jNWmJZyPY6iNMUoR93xLqMwcv+E8X7Xg1+Qe5Lw+xTgjy
5OdfR5c+nMDiEZA4PO4tvnbj5x/+SMS1I5wrxNaMeqwd44LGfzmVyKfiSLhsj2eJ
9ReixsJJ2EzfYJl4BkYFOOfTNZCcUU8U/e+LzXYQjk4EPncaFaZymBBojG55IUVZ
6ya4NUtyYqTafqamJVoyO/Kv+eXJYQXqSOHzy+vm9YLRHX25oQA65quOslyCPK0F
fp3XELKeJ1vLxeaQEghiQmnU14CcB7cV5ScKfP12xNMGhUBviabINMkGWf2M35qu
8GPrOfenhBCfTVqSq+A8guOLjsIoLq2QRZkK7BLxHx9PNfMNkwMJUxFIKPff5tNB
P5O7SiqXSvp6w05Qfr6g35USQLSebD22VpP9tFBjwVOKXUerhQSA/ZwY9GZ5SXEk
49i61Q4lKafRGx+XxZ6ck1yzV2LaGE5X4VTxOdqAHWu9XpxxzE/QEydc+fciJuo4
j0rxjIFyf5KiKvh9k2n4sLvEzkmwWkL4RwAfLdYGmkUGrc83L0msCd/s1a8wCVFk
44nIJGdWFpXwZzqP4Wc4gaRppL/bAHKFuIo99msUESTX7Q9GGf78ZXewyYg16a6U
ymL5oK95SYknoyw1mSGhupNrBJ+sPS91Jr4+MZ1rSJ7RyrkAZW0V5n0VRIOCAiTw
gQ0I4ZeNceiLE5SBajkyFBd72ssrL25S7ta+cYJ/qKZ7MTnMc4XsIusS7Lqq1xq/
bhHNQ7SGQrGE6++aPxaXJo9v0eiQ6lNBOSphGM6rsps59Tr4a99O5LgXflCNcitj
qwLLNnL+YorV7dcz21bK0yu4WWaGYS5RREVpTbGNxhcbqNjnh8GfUg1SOFgZnefM
Jm3nz/XH2Ra2DeBj5EXO6GEMA8FLStDHr+tJI7r7tQrh8kOEFc9VqnucWwJX58dL
OOugd0nscqIl6O6iPdLYu5tJboTEtp8kDZpL6BneYO3NoAJY2G1wNwRrR1mrz4LI
/boAJ5/W6QLzqIdrXIRfpXiRw61Relidmn7jx7fEC6CxA6OzqslDKjDTiAgyXu6i
Lqratqr+ev3CJYPIYirSKo4Hfbfyq+1oyzLuvcuW88VgckdU2bR+n19vzjL48GkS
HPfL61v6KTjQ64xcyLiXe8U1RpetVERbfRc8GA4/wbAW6MZczNUyeMPeSPI0/pcR
X9gmaM53Lk/LeLpVindd2oHWn+b8n3ntu3msCOXDeUZDm4MYhEd4M6N98o2UOUVN
nbTjTMW7yS5uR0savhB4k2pmGL3EFn3KSRc79/dur1PzZdcFx5E0oo1aLJcmGlD1
V79SF5KP/6ssMzGieoXab/FOfRTVcgGPoM52u9tpgFWHHdXGHU7PQFj6U6TTUShF
mudqcn96yJ5skIGSmwG/wCsy4/mNH1TG0BVto1saStidU1B5vSSP9wgUjzs6bDFT
FyPZ54roASrL3Yq3LziveChmQi0j5YTwVWknFjEdDpgyZcwJqPUgy9HHXPnly4Wb
A3NMydQBioWgXOs4Us3MMRjuCXehdYT/ztzNv+SQcSut7xfCkSgCuELn3EX3UmIs
rEPweS0GU02G8YCblAjAFhLv6pXpLRjInNvJl0Yhj0W2EGdUTz6v4j7hwHjmeEtf
5JzMV5ccG+5/Efvxc4ybIW/5/nrTtpLTPZ1GkOYbU+4T+32pwjWJcsE38dxx5yn2
cxAXPsTAfxh+453Tqgbdz23x7k0LOrq8xGi1JWTasl98xrxcgjJtbX4GfWkAB2DT
V99/SapP5/rXTezrH+QxtXXi3ZUKU+YxOOhmPZMIGK1rtDSXNaN4843TFYNi/Rp4
QOx2wVDA1SpCVzCFdLlLDzGVvIW1Y9chS8QlxxbQHVtmZZcKSZbgu9u6lM+pgP34
aeM1lohaQGqy/K8CXZxig4hCa4EdTyTQJ0VxnodVoOGUYG6Ydty1bf6AzbCMue2I
HeVcTjKWOY+h2A+WQFmDStNLGPC6PRmr9tssIfWnp16wbe9IF/XT9XxUWczX/5Zn
RzPrZMbQVS3NjIC2mo7RFXZqUKH1kW5o4lfeSd8jj1+hv0/gk41ZyCnTXGWYkmeu
z7ItCtPM6oeLUxOCpqoKpw1MkK+PagJ25ayuWeZ+rP81ghwhEcujsLpxBPLC9a7c
FGIKT3SBAFo+WgHlvht8JK58ntL1smfDtwfxThdvkdODVPjn0AbhRuy20kHwC5jb
g+IZ746SbEpNSRrj/ba6aGbAEgtpL9bPJMKZGz1J2OZ9VfJuL64xqWF6b/ZUKWvp
NXltJnXSeUbUUedtp+uuXCif0rcB0KFD0Y8zMosyKXX/fgywu66bbKdyF8jqFkgJ
Ma4qVDI8/kYY3XhlbuVQNCajQCNYm9WyxhktcbPvmfTdCEKTDRZzQ7OFp2BLu8dv
HaKMr8PGb7+x9Ib0iR12lSSEMNSeawpAYq91PFFt+TpXG+d1XDaE5LUwtepJELVN
ErDfS2VNx7MCEkpMH4wKWkTNImaS7QVHMzp5Cwty5POCAc+1yDeVGjJuOQC+NrkG
PLK0kstVnj0/4rkRFfeKahhxSXXUsqhF9fAhDcMOYp2HPjBbZBAKqnGiFzPDJDtG
9b7Asd1oNB6qvtAgtqa0IGcgnnNTyF0AxJd9yyuvlaPRhEYXcLBymg5NFpzv3WhS
qUoFzJCU0+b2OKhH/wsCVzF/rvF25T9n5bEwGT1QKzvdViMcYCBSJInNZDdEhiQd
DJqCMDeDQiUjngWKW+eNHKWkwnB8fXzx/LZY7ax/PSu7acBcRrXMHMNocDbAt/3F
KH5uLfSQ6PPCoUD7I0GI7AB30ByGkz9n7IPh8dy5PTRwFU6gL7BUhTOeowrdcZCK
GOakKLAwGOMOPCP/ZT8nPWPIZznBZMAv07Ddsb/3xkrbfszFABg9866jag7NPUdd
EOUK5B0sDm20OXj06/2G3K8tD3pmkpT9DHaqigRWavZVFOhqrO3K0gx/ctEGoTeC
6CGw5SMfMXZsOYQpyOTFcToo7QHXIWx6/VEQQUgXLacJjNeFwXkemxwtZotHuo6k
VWYzwZ1Fh5qI5MaA0ob083W6aLR9VTNQiP6UAq8nDWxi+nuDI8QhZv8iq2cKx8SX
A3e4Q3+MhP4c89ASe3D7dsZ5jv9ev8Juo83nvnaPs05ZHE+J2KSt0xiguheU5GtK
8gfy/RWQRc6MvR9mbmgWquFtJFXMObimxOEJGhttO8pfThA7lU7YnKAblJvCtpNc
FXbQOyvfhm2KnLundfungNrEbe1fAhMVvthkJrU4j29xWZXOG7d2z/LFJrC4OGKs
Sr8hCmsRI1jikT1bp5tZA2wwQhZAjTw1b+SPUsVGLkuEGQgwxNog6shvZQlnXFoS
hQi/PxWfaBfeoQavU2odh529Ab2BO8ijnI1kjuNmWa2b5y9Q1Omw8G8DIxnW3Cgv
8LVvHaH309D1DiTqICYfWruKuXtohvhEwdbkDxceh8htmCm4hGlvhC7TR46gk6Fq
I5HYfUTb46GShJHysWZP/W1kz+pkFkuwAzSlBWryFHtbTrfAimfDS2eYhcHRZbxo
rjzXLNvJrsxEQok6y/JkJTcF/kUWAjA+xgOjyYLTYCClHCO2FE94JuYX9yMLxi/g
eBhJ1/oFDoy+9Ghk+DgnmS3XIR0YizDZiTFHsnlfyV2TgHlK6Nx7k0+MSoENZ1X1
WxPUv3lC3CJiHh8Cxe5rggXCrYfjaeyT8MipfeNuakel25SFNXryYWDdp8uIBSbc
p0A64LP8ejlhSAOcTI0aOQOb5cnGwRo1MX+suNPNCHMk1gKqfV6ZOloNC79NvsZm
rh2/K8aIMG42FJJ2DaXiYoCnJ8R8BozwQjauQoqqwT9uwzhcUWPfn+VeO3fANL1U
8XPEjM6V7wHPqhOlH5SSpNZfHQEe/VaH/rbMNd19coz7sqpasqsOECjxjBAEKBIL
Vjvli5gRq8D80z27c183gOP9kVQd0sOm6osNyMnFKn033VPZOYK+un5YuCUKBMpC
352bCCm/6oMibfRU6YtYsKBXF7bL80M1Odp4dQISrWI/vdGXNpsrNRCPHwkKq9Zo
XFHL+UHVP10BMDOevNFOVGwfp60AZKOtHBAs36AKyRM50HinqBU4GyjxF2W/w8t6
sCLf++b4O6CIHZU4kmAI2DeDPjMZU9HwMJzofPI0aTDqlAN+xDrCvom/IeHnb0WA
9t7Gd4ufybMtwkYBYNcPgjjpOBnUn62v8EvhaV3yJF5YHZGSLs0JoyUELN9AkwM5
CeEPOfM4lmD0MuXRGkSTyWhKjuYe79joakB+VWdJJo7EkPuprdhNtlTjROgMZRN1
dFuh/rQht1fbB/EhdYiQb3ykhfWKvGEwmv8y7SNO7AwNEAxlhvAcwipxOo7F3ZGs
STs6pktfzAGwruZQAAgyMBaFWXYriumxYgqMsTQzxcfMHY0D1efRCldUXr+p/l1P
HBnPsBqfriHB8zyiu5yt8Qe1iWLDKaJJSTORsdV7vN+iSTJVx6YVfAKkrQ2Z+ytZ
RqQmRAVA27RgdOBRQ54oSrdDMpl64oSF5ZXGTVO7jirU2ykdHSuM3fLPXrW07byl
aGBxFAYE3Mmor+bY99QpJeQewpTylYQZW9vJi/q63CvNuFs8ev9RqT1lQ1NNXcpt
/KfLzBAr1r2k/U1tu9l8MJrJq7XZyG/WAdqVfEDFtXC2HvhK+0bN8wsnbOfnhv0b
8zeohHgPmvSdLP4oe7bhrGjv2ci+Gh3A3JIDAud2ghoesrUSuyGCuR1bloStsoJV
X1+NVIrjDKfa87w8uKyOXJEOiv18Dl7VrfwCssS7tTsHvitMbnm8+Sks4rmctQOJ
uez8VTrEFZB2VGHhQaco2SoONApBJpf1EGhjJg5OOvj9bax8E5gnF7rgiOLdsT0w
8aRdUomAkAa8W+HdEypyimVtEJHOLrn0QYEIvCRqmkxhSFKx8oyAKwnJzuoIuliI
D1qIWBXKCL9JWzjpiBBwnMcRbu5HnXu9KHSIcvvZg+pzyNpNiQDvTv304Y6pBLJA
iP7yZOKOKrI6KA+P3ssJdxTfscvABAGTHrVqrI61vwMh7I6rA12Aym8rm+5C9gq0
o86o+OWde9kHW0EYNKg2G/UFelYFezf5Ej7FW6hMoeJLTyX2BQnVejKXe6w1b2f9
gzl+hfgbvyL95q6d1kytnGE2w95N6ZAy6SuFAcLRRRY1G3DH9CFKwKdQQJftXhe6
EIv1qm9JS+67oTaAKwQ/Fw8CX/7URs6IoIlgbXeACgwD4AiHNnOz6+iBTG5/Rtzq
03MLBrwjyPjZXT1ou97CyJqxGnYu9PFSpEG89zr5J2JiimGJHamjBz1gXLLyDx2H
y8IbDBHx2Luoj3MU5xzPTIaXomWo0DnWNME+mQGsiRqGuq0GaiProyzVZiOkr5Ii
oETm7ben7KzBJf4jPEkL/fgOlCWfZTK5UXynfCbtr5KE7Egeb82u2Z5z0Dofful1
l2vlUWg1k1/2Rq7hiOR7Iw+heE95vOccUMBatB4YQy05NrtHxEkTycXkfhvuVaJ0
WNNAXiLvcQe1s9tsrlK9YHY8ELwHlZ9Ofvxf8QLmFL4YJyrKLhWddKe7/OJC4JUb
xVJTBFXD5NCERf9usGPskYM+sePzCoiCA3E1QHb0rA/JMAnjgA5IEwIOx/KoIdNm
mOG+za0siSpS7D6P005x0vaLfRjSblIUUtahnW+tOXE0hn3TwwBcdAGo2a/3rYjv
kUYE4kSwPbA2jsvF8V+5UxJweuUq3PMdy3azDP6zLYZAJOR4IvkcmdFY473xvomz
57soXZQO2ZxzCpbuhcIs00Mk2VL1HOYXZhfXJ91R7NM357nCShof6vbKqztuNNjz
oKQJCp3luj0XOqw4B8WIiB68b+ywt1XFrY+qyKwIr4ztTo7wkFDJ5tYO/UJnpAfi
xDQFlHI7qu6SUF57O4Ne9/Ul5klvoSqATKICUK8K+2HwncED+A44ZkqfM/kAz+DB
tmTW5uUUiumuoYcovM/xQdifuwMeLabaVXv6VL7oOtOwZ9UEIXfwmChNrECb5QTt
QVH8uvVtqXKuAOvnnJ+c2/FZEfqyuxUpzwXS65bXoQn/QzPvUHzO4yrRhrHpLa3L
W+dqAGu/M7d0kVIuhHYr1LTt6HBb+EjRLHzegDnxQGv9WGhv1AYxjSvA29ogHm9S
qi7OTpGpmN4TRhL/rU4jyotLmoeJ9odb3RPG7Onl1zawyTiRvbCqY5u1qj5hw0Ra
XMCNmlPahc8A6Er9VgrQYRpEtCgnKVsBzfVD0B/gCEvllgLIPxW80mNdPjMayGEN
rg+lIdpvdSgc5T2Th6+zS0PdZb7IwKrbbDa5TyzFNTppS83FPN0oAdTTvPFF4p1Z
d3sH8I4bWHswEoJh6cmFIgg99anrzeLEzECu3UhmEaeKkAhnI+D8E7266r6wnCCx
gVKxdujNrUvyXmRhyC08nL4qQTNy5ksSTXFuoG+X0vYw+5/Kmthdka35tiqPqOXE
NA/B9EPhdDk/wE8+4gIdcn9yG8n4AMjAmpj7wWOgYmeMxR8g5r6efSGr7mOPTHFv
iE1BVB9K88Gge1jhMG2mIv7aGqs6r58XkUS3kYsGiPvc4uGDV169p62zqHaM+ZBG
tYl7cHAceLfRBcR9THfU+t57JjfGwB9xQnxnfctW+yQNoGym3Bm4+HDd8zA0tFqK
0SNVDwAoKI1C3I+FN96yW/KD7zGc0JnUlIfBJ6LfyYwDfcx5ek8ibtJO0XWCuhGO
M17QZfTWBRd7lbiU1NpfTbuRIcTGk+Kv8wDqgad9LUtVKuhR9uLAUbUHRS8Y+KEo
QHLK3dCPiOI5QSRrADGdpf+i1XRSmVwmlmaT0tYpGa2l36X+vRIijlyRlb8hJMH7
9fcPrP2lAQ+73bPfTrGhfvc141AhppGlOH4HoZ8HTTOiLIZYKbHuPXE+5u/lKoaZ
TPNhomQjVmVanyNW/CPA+g/InJdyzUgXs5U7Q91NiiKu1qz7A0PM1kpmTtaN9J3R
PadWKBEnmNpBkxlIaEaCEqVkl8/jFxg5FR9L+QZJZhjcfmy52NmG84kwv1YIQMtg
xkVR79XIt80LGfR7LCrVc674nXRlBBcwnG+/61TGDsyrZsH7t7Pyo8DTQ34yhjp8
g9wXk6rEZ2O2ERmzhcTQ/nHSABeZZVpK8QXW2Ibj0fXOAtJ1mpZjpWJeRJCiQ/KG
QkvFo6Bd8LfXRlnGK5sLs2tau2HgDN6nrF4Idj1VSWMyia8ep+15QCP3dlPqOQI3
GF8uMJH4nXbCpoX2XW/eR1CHYCi/m//WwEvgiy32JjNkp7Hry3FMzbS6KM6FY9Kl
dtbZgAikPpWCxGrxxZKd+275cZ5OV2VEzaUCQwD0IdXwZm+DUAZd2xVw+BvGdJhZ
ZDeZ4G173ApWPw2n3fjU685iyqlnYg528qPVR7i1p9IwkFrxqhZkHx5o3KSRIZ5y
ORB+TptOmL2D6y/rsrDca7DtOuoAAluB5oY/PceiRM/zrcmLIzbR7Nlv8xZOHhFG
4GNcXvEMwpWAInLjfb7Sgi+3HIUyt0oBX+WEncUVwz6GW+dRO/zY5JhlgqcC326a
KtIpBvPMT6r1o4WPTne2wOuQpNGgk8diwOJr6dWWOs140Vq+/lsmRqwHBbLzMEml
O/7g/rM5LpSYQkWKz4g6xhlBQrC+0i5mS59dLGcQSOFndjVCiyGwg4ZF1dDfIXn/
mWtOhX+KFSn6jm1xm29zYYRy+9kwGV95TC1YsgS+rAFAg9GR0WUg5HL1DEE9dyvf
V+MbjCYtg1V2ttCQCfo+JGCqONHIiHdhpm5iWn+uEDu86zNexMB+UHovmwG/qSOB
f3YtBLN94GWxGUiHXriInnH7rrIhqygXgpJnjSXeuhn2eMa6zd7ZRohjBvrDuv3Y
oR5jEAWV5uU/0eklsK4hnvJwCTVa/yXgO85eUvmaUfqOtZ+oJSIc87iJHnex3qbg
W3nCV9fYDUy2NauosJUCZ2LEURK9dot1Dfp9YEZJ4fZQRiDFDXUPb7tVdRfkYuTk
CAFSXe1/qV1sTbE3kLhBNuTyOlI1bHSCnZzZ9POlZuEQSkHo4mGi9vncq+cJb9q5
oqOdV6DABhx9Yu3Xgp8pzWn5b5cXPyIDfcbym3n3/FpNRnrYCMQ2/WmdlSk3StZ3
OBs3/WQaoQ3Sc3bs+BE/sxwm9gCiN044/xu7Pe7PPeCC5yG6kDtJ93DUavxartYK
FHrxlzNcOAnwWqpQ2+fX3/DO6Erdu4bffBvNiA/Vwq2fY+SrejQvwz89lNOitJQK
aU8n6ofYCguK/9iA3SJFAHNTvxkKOfdUsoIUwijbi2RAMm9PzbbF6+NqP5GS/2Ck
oQ3LE/G7N8UTiw4YAfU9LXQj6ZiwL53lPGtg+xUo1ofWedqMLyRHTEhJ+2gaCUbq
sk7ELH8kS6ePMxKLbMBKNZ+GCJ3SdExBcvfX2Fb5lS6QoLGVaNzrGI0Z3Qva/8yG
DS4k8X6GtYf87uLE3bK37BMwn7Um7F7MaNlxortbnw6BH42K62R3HWjilHH2JcPQ
0whmRFsAA1+Ea7cFNADt22zfbHEBij7n0CpxHWPo+gGRmRrTepsbocopn0xxVB2H
POJozlJHhDptG6rqByp7r2EJDaFgNriiUMQHCkeVJ7miBwQ4OXxGGvHrPTynLKAl
Dg1rmnM6oxOVK5Cjqh6o+B24nhI/6a0Mx9oN10r2t6R4ZKL7NFiJfLvd7BIpn66S
UFJq4WOaWGcRKoPlbU6Dw6kdjWdAVLFfpkanroGwch76cEZTXtxCilbBLhMMZQaQ
RDpDcYoyI87FqSmdG6J2bTpEaPrRxBXWtYT84qN8/xmpWjQR0Lljw6qLLJCtYKBO
AA0Lv58dtkpAGiTCsrOxpVnFzPbTnxeWgsogreTV5uzwyCWf5mTBuyUm5ruVMtJG
0WpNBk3FT+U8wvNj4QRys8JTQGF9/wifT1XIBXZ7FZGyhPzZh4cYzR9jT9wSybwq
gqYXHkSiucicdaR0eJwJF7yDEzhMyeoNuWPKWBscpek5TiAivaiLmRPzQhSS4sz3
7jNUdPQGf065xI3HmUhK/cJgt3dFzQ7hS+9wjeluW7Ctx5qcv7F59dnAc4Ab4s5/
bMZ3zuUmYC77U1G1WVblBP0I4uEOPI1cBMXSg5ejRt/p32wo+DxA4m+g6lSYi+W0
4ln6eOexPOPvmlHvqSO+x4+AzZRSgCM6mPk4mLT176sZ8UwrVZfihO7x9aDTTwIn
NWeOKVEzv1GllbSS25hk5PtesrzWcrW8Jgs+xY6KOUMW1uMV54nBD0ZBqeo1P6E2
3ZLwAWgBU4FRBlfS/v82wsY7WMo0S1SF1jGFMo1DhkgXRx/e25fnkBZaYmN7rNA5
0ehpfhhefLe0YAPQKLdx+SnJrzLYZI4T6nGzsKjYKchdxeA3zyYEHq1IbeahakoX
Wkhp7NtgNOhioGXve6q2CbtrjZFACA/v4GoOnQpPMIMhPPKvnd6+Wk1r3Capc4MA
dCdrsRBTXHh0IK/kCCyEoMIQmOhFYMIyLlTUdhXS7ocbTZECfi9P7Liom+RsKJDz
+VrAXv5l3RSBh9yfICUuE8+oNg8l3+sB1roSPfj9zpb0x05HrSLLCuNtwO/YWM89
VjZSdDvejVfiON2Zsk7iVwxRLC1e/L7Xyp9/Ss6BQ4GFdP0CTsLBqIhfTb23BgoF
Glnbn0IwZAblzdIlGW6ZbkPQayk8H5eTDIRyV2gf9WT3FAfJUUnXkcNlcNU64Nxa
pW0C5wZp1D8FSoII4OpsAO7Y6itHM10idEJuAgcJfWW/G1lZMcJzV9Z2MDMNjbfu
FWw5IU3DCsqrDHq/gAY+WLIq6LP9XF93OJUHjc/u/kv5jo8cBIkJ2qL+lgEqY+pY
kni+PdT+TutJTR4jQwuDNm3I+OF0tiFbkGcvCwQaYww7vRnRKwYBcWwfZ8Int03s
1LQM+qtE8RT7X7C6qk+aAcolZZa8mJ9XsCzFm4DXFYxGBc6FXQ6bfJsM9YCjJuO2
PIoA6WV9SriUXbtkMgG2NMxUlU7hkFODlVNFz3M5EPTUx/l+ZAiJCPsKzlYuHCum
D9DZGDrA5hvwJeCbmJWqIfPOzYGXBEuiTFT11fXpdEKFtE0Xw7BdMCyuSj5roG5Y
VHrMa6cypTv5j+gZubiZrV4H0zh09bcbMB6bImX8cMavSKRgf6k+iyHtcrfaDUTk
685zzvEniDpeqdLRQOcB/BydTRPAe5HMZAr8zMyT4hh+L8WstHkmSQ/JWZmKynsu
LO8k3efq1rSW04/Wy5nYCBHNRbvmMEFcqKBjRqgio2QG2z3stIKg6HDBneySAQmF
87ehk0FgankNhuuY9qJkFcMOirXgKKlTmolkwwHpWl//pDS6mlvb8P9KcjUlSwku
HiwXftkTuwKOk0/A50YD081JUZgOcl/V2CKlbkdXSNwUzbfoVbXG1TiXgtGslrVD
Ugih2NkHxkiyKemD4xQ8aoCJG+HJUX6kMv+jruKGrwPXGkz5j5zPw/UvPtB7s3rW
NGimVrOf6UmD3S3TnCB1Fih+acvA+/GnI9ZpPpCoESrXffWtqiWu48zI2LiHpaCW
zoTjMYBVPPuKOAY5TZhB048ePeVHGTUti+wZA9V4pTssOphIbyYsq4ZWUHiFALcv
rwmY/oSxFdvJxcwRIbMnpIkXM1v+K+e/6AKtNrgKtTRp16Ff1VyNEPW5toRyuGZA
fhudpDt5I2HfNfwXBNkZAfdb24F660ReYAYKXp7G2yr6v9cRXlCERcj3pjy2NWeM
sGOuCrUIS2IS+2UYit1tChpYaAz5a5Ij5L+ydMD8l5Xu0H76eXW+acFmo8Y1+mir
kMfBm0w1VIQV2d/eCyLXJpEncwiMDu9ahxvYuOEni5YunpZh767Lc+wfl248j/VY
z+3/DXuHj8HLbVxIWJHLPiPs+E7N30XYArWEDI5qmYTZIGpuvVHbq39q3wPXpYAM
EOI7B+cijFafhoyn8rjZm0JLv2RW+haqzVSLErz8P2qW0S3fEcVLENCyS65CAZjC
0YqJmv9npzFdqmyQw5bJPK2tptA56KZG/yDD0FvmbCZZT4ARNRz4aNV3DAt9+QWi
afUC/6lmhso3kL5Wz/jZuJkBpAwpXz//hv4kocUuPdwGTozS+oO/WuOC/Xc0omHU
TygQAHis7O3JkGT9QaaMLp4QyC4HcfHpwdZw/1F6LumoW8sVtzIIzsdVbD1yrPmB
pgqWK5AB2kmDRglsKt2iFiIcaQzt9uGJQNPcIWfuikNwpbKm9oht+D1j0m5W9u2v
/PswyTsq4AHARVyQO3KL550FfUOOVHPF8nEEAGSudDekwN83Sudw+PehXD0ixZ8C
AtawGTJqZ7USqY4aylc8ZgC0aRjPgu73tuDssPqNSWd9fmYPvU2bJpe8ETfr6+aL
9WOnCgkyYO7AflLX1R/bsYOR4qxVQrkYB+tA1Zgqfvn/BJm3XEHxUzm3fQGbqYXq
cMJ8OCpMdDmo5WnFlslqcp4cq0E4WkBWekmk1ngXKPVXd7+tYWpkEpjfPJTLmnnz
UBi/chVjz8bSUU2MkRKLsbUQ3VixYmKxvW1k2AfY47XSkpcGSrfbJSGI3oaPUP/T
4JVBPKkNovnFQtk7MayBciMrdPsRyANFuGWOb13Yp26zSUqt/QnHskYPKlZ4uD7H
FMJIkXvJ0oHc+GpcmreiGSDACvaFiBkPVb9jzXfW6wvnDSRLSbAIWBSJlE8+kEus
zQdFiCYW39LWRpRFw7ln+OMxTlDtTSvjGJydOMjD84FssfNOt7K1GTWmB7WJ6N8K
7KhbI6Je+Qk3BYZSK62gisN+H74Bavwu+Ei6E+IYLw6T5o+GHX4d6cnBW3Zhe+Yz
wPC5vrBs6f0F9yUmNSe6pgTwizWl3R7O0HzJGrb0FW6+8QHS9L2rpxJV8V/WZCBz
5+eQzOJJxRUhBvL14JndTdVgHRoOswyQvkEXeit2hOQ47r7IGpuqVDY8AKlO0Dpp
I4lLAL6kdS1tcfOaQUku+uXFqtYxfiwcwMJOdYU6VdvRagoSRmXCbHf7yWkVSELo
ykLXDAg74A+7A76o8rz3XPGpusFxTizg/iwtzci/0EXKAcYzSkZZrKXqCljZdmfw
TRrqJOY+rU8gvMbcm0XJZu0wZ8NJkY2UY+loiyFHEbQje2l79n7MZiBv8lcpIMnh
YLh6OfPDkqcsUWJt2SQv+M2lbaVFIVAJ2JLhIziq844a/lukirsYuVbHEaJ16jZV
FBDeNpGTqq3aatSzYApFkG5ueBB1svl0PYGAoO4WK6vRgLixODTwYYaXEtFCRXCj
qIpjtQm8qYC2iX3ZDE/a/leETI6x3UcAf4HGnknxiZl/FMNDAgARj0oLo6wNdIJK
8yQWZ15o3QFD5rlE57Vti118athX0vkhiYtyK+qeJanR68Bo5WlmxNYToQ+MyfRJ
w0U2zlYTPUP1r2A8wyOSaApVQi6norXUZ0kshhcdOycNoBDuAFvheNKABx7U1CCR
o2EMcVJTzKvOCOkVSMnfS4GAYLiB9Zsr4cruDFdTmNaWDfWrK5BVO4s1M7WkRCwI
CSwfO1lt/5A/Ffz63W88i5BOX+zYSTHAeDPe6eY/wRh8scS4RMZy8YU6J02XBruO
APEaYosJYRovAg4bLoJ3KHidu1lTUdu2eVAGSKokXt7Q5KnTGHDwBzChdu23ugs3
HbuV2n/dwnAlTfYVlotWly2AXq1DVkJZ+pQ7pNAmq4X4EWQnh9Bh3U9/3xsXx9JK
fzuik/3tfEYExgi02SZNANZvKEVD4DYJ+1+o9h8dIXQjTVjiSCywVXL/5PtjRS1c
XljKiEgBEveQs/Lgx4dhGYdkhXW8snODaqbOUyVAGA0W7661Kfje9jYoqaHGybLq
o6PKi/fnBC5nK0UIGBTLbmjnH91015VT+NSygfWOVNhnns6Xe0VuUo4moa6ThA8+
duYoCUBFvOUCL/hiFgV9IKi2jWg3ehRp0I4na3sivnVEGHpUfIjGj1k3u8q0j5Kt
xEiCn4rUzvsUMBqN+3ohGfgazzW2IqvHnFbLHptph2biCBjd81yOrf3JLN7LHEDi
TaJ9h5gI3amkNtHI0FoAeF+4SjxFqgCdRK4m8B5kQU5u+0WHbU56OmEdfU6eJ1ix
5GLtHK/IxOIpWzqH4sUlP0hbq/+IbVG1hIf084cEkAB0R2TVlELy4+gBh3Otueth
baIDXsI8BhdQd0+8SCR+UQvN4KcR3yvPue9KBu7C6aeYWQSydKHaEoZ3T9zRb1Bf
qqaFaeZfvHVTdGPc1sFgVU4V32MUI8ZBMUTG4B61ahaXuoXfv4tB2hMq9vm2lV/T
s2BOgBPYnSHSjoUfBQWPPtyJVRFlTkl8feAtZxCpvLAoR8m0n0UeEpTumS3JQdF9
dJREy6a4FgeIEQWg4pF9/7p8VndwYPwi0lEeH5MoOFGBazqJK3EpIrA1Ff2w6DZ/
YH+fKg0ERznoFquuye5jEy5cqqZANUfShmKM9h1J16sg7eHRmI22VUzXx9We3cFb
fFRSXtcflt9GBRFGUXn6GESxNxg42LXuBaOxonUJ+05wzfjjygZnqk2wNltaPnh2
xmkN+4CxECtXTHcNhTwvQdXOKx/z7jqrkZtFxktUBJT08u+2IgjORpbXg+obNWX/
GGvXgbakbxuYL8dCjtatW96ZtJV9Solmeex6k3fppB+PFPWMoO6cgdY3Kl0nApFl
6D12kVGA9/8dQ19meJjTmrPDajuhZ8foATf6wwO0rCXItouWIl8hJI5h9Hr0ILmu
muH+2lK0q69Lkol7Cc+4TH+76Et8r+wDJRlFAAlBUx6Wwcua/mR89OxltCbiAH2M
HKyQ+rcllXIkEXz8fW50+VdRWzdydvhOyjybGYptCrAInGkuuJwypdo/e9BU33+H
S6rcNz3M7g8G8kAWNb92ATcbMxHkyNAVXq4Imu5vFPvcXI+QXL8O2ck/BsFp50Nc
H//WJR9sYE7YYKAfMxndeBEXocpI7nwPAst37MI9Xujia3pCXViXTgnWBgRqfttv
E+jIdTl2IqlryLRC+MzFsDBQSYMDJJNC33lnPklIJwTBK+Ss16x4BTAlZ8pn+MDe
gEGTsZBAEr5pmH4WBgmH83W9KGRh3h708Ta0M5pNFUCBu2nPSA4PUL/dKtXXJmAq
KOHqrbqDpqxL4vpXPunzokmaT332wwSoHZiLvwfe4dVrY9lQbsj6wg89r1jA3kFs
2UHpv3q0m0sIdVu7joWa2fwNC9FpeI22ZDBkzQxvlqusanWrTNkEK0LecwIN8iiM
ueo136O/4Ln1XS/Qq9smVwr5ZWCiQ2psv/5UJc+FdWltuvtUkETzw3OiDWEx7ZVE
6c5iv0wjEuAi3oGKcFHoQfWacM45WLlnUOlRy/VRaK2Mjys2XKoRqWAivjmlgbn/
SaJyoT35b+Aj1+j5XbLs93ex1kZYYuBDXjK9keWk2vn0VqCY/hzLAJQS/blAGNUU
kjzBeQ7EC9nNZngJL7VmXfpxutScRzUhYmknMxUEHToXg+GNJ8ySs7BKwPmTJI4L
1IuMSEtGig70+dQwngMn6Vma6+KI/O5C3BERPW4O3qLCOgMb4sRALjT/qTkWlcK3
vy+kuKi3hr4TA2TwErVWhjLGu58L51ijKrD1vq+BR7VawvULbByh/6NTCvID9yv/
nDjHfLRsWhJcg6sSTxOg0Q/6YLk3HXR4LYJCvTMWDtgzmyuhcp0B6h9PKUJUZB/p
ByyT1kl1seOi5X6Sz0WzgpBQskqvkW4TY0fUhfBerY37doAP2UMb9X3qsnUe28TK
fVptVI6G4kkzdCcV3wkCuKKPA079le/sEWr9ckl27l5q9fl8tgwQrA+dT8B3v61H
E6rxtN9mP+ht6xcZFfndy0lb4FOg7FYAZSiYS4HdryS3mhS//kYpxP5xXXrKiegK
I9D+yXi91ENP2ziOhfPlinByTDoMvuS3ONHW4erf4w2jSyYbIBWHfxTC0FgGtwh1
IkkVwMxT3qU9GxEPVXPhO4Ia9RbcTEXVlETh2mluHCjf2NwxA6nY6xxULIA1f84H
q/AYu2x1H194tkDnVW5XwcaZC2rnpLUs3IF3g5Sas/EDOmyiJuf3e2IRGxEHdLKk
LlGfmkVUqJ1zGT1h4RcelqvirlXnqZcvlqLOvRaac+/DYP1ZutV2fPUUp9i4hstE
TS4fOvi0xIm32t516pIdfdhbTJzSRYDDxE5sUgBBm1L1MxbiX5SwBOWNHD6RhM0+
9fBA31UDRcIFREycRtD0a401ilRmsT/eOLFSliexj8Hde3IM+yGSa/eMiSsYkVpm
5QxtuesUCmbAFZ1Es2d96XDMfyaLoMtmuu7f6zFap7ZNGMthJ0MxGtM8/sDK9s+s
1LdklyWc0ptu4mHICGH1gh0kGnXx0unZfD5Q9quDw7ai8DYPmjFnOJBFKa6pY7UK
VdgFfzLmukEMBItrm7EdarPIB0hyJy2Tvy2NOmRuzZs3VkOk/gPqu6y4GrngL3QI
yltAffQZHwPHXO57AYDN1UdOFKOnj4B0o1Ds4dhNv+AwrC3RZhERZeWjmPkn0xHg
hKtT/GLbGLnbUxkSy9AYHFV9R+ftzB8slvzuXhgW/2YqQD4nr7gGzAmN2a7+x8Yn
xdTXgDJYZs8HtSeN8sP97JIAYQB/ykjuJfLL6k/IfEH+SzrSxtTA5CjD57YqpCab
uRVTQMChtjxZP1JMK/h3j72La3E5g46Ap2yLe68HQgApERF1PbJaXzpLvEY6MXZ7
EX+xF1Y2jXbgb7P1NcoxUt9+w+EvpOlNL4n66Z6XrzOp6wgRzV/Ox2980sHpBgRB
hx0JTa0lginSbCy9JdDAx2ISLAb+cW/SWJs1iUEsLKxAkUikiEIQcSchYnrXNbIW
UG/m0GUGT9RfMzxvONj1GamxCZxnJF7cmVCi882oHdr5zSdA9eqSLMC9TTxqpIZP
aLuBphyeKfMwqUqcaB6eNEBY569vBZgYv8CZ8wna8mds0nDevh2vurfvlbR/OD8Q
7BsUg46CamAZci03eGzkk7iH9FfyuphlvhYXmCgUbjCVcNLtVpmXrVyo/8eVpxiq
WQNntIOfHAIk/LZmnUIsq4yDOCO1W/KttaMnxDtf6St2uZe6ctlZfaj0fY7cvbR/
YesXHV5ZiI2LNnzpS7WrwXH/SRP0EolkG9O2kmbroonCwO2pCuJlICagFR1j5jvX
8sD/J8RBctArYo9aifG3lkzxg8hEc5E7+nUFUYwXzzt9rFwo1b4Fzb8/pvR5XP0n
Ib4zM3y1VdQo6SRWWucMrI/VCrHxhpxLk1hc81FjlQfWEArvEr4nEYwzn6ZK76aJ
UAm22ekVZZRceJH6H44WgQfdeGmVQpaOwvL69JdEUICYBRNrJQmW8en8J6CKQEDt
OYePImfHIAyVGW6XErUbori6Kzfz2UPk+gDUrgDn/3fQewvlN1jHI5DecyVLIrRl
MxCQBdoU4ck6RTl+/+b/r4JPkwRiKjXg/s9AJEAL69nqnf2hPxZ0I1tQOrf3bvCF
r5ANm7kZTXoPmLsrHFYv1IvQKUWpxwym6VxQKKNNQgfjEAmqoMpePnvFB8t7tzOp
AVpedCOWYjfBO+Rl29Nswcg9sCo0afyV3RR3bwNi1lgk4SwlVQwMul+ma6xsc4A9
hxa7YLI+gss7ZRZAsNY5XgE+Rvly9FMxkjgWq3tQR9+AHYHRAAPNOzy1x7HxP5/8
9m74wjasstjrbq/oxi9CPNfSWWV2TIVk5aNET2I6lPLbWwnj8PDfPSLyYFB6lkWO
POj9T90vF+8B6LCbVqJxTqJMnj8gw/T8lDpCE3TxaZO5Sh0yGWNAFPy/Sw9OWCNb
nVLKL3bqc6NSlPQiqIht813dtBlv/MBJZOXas8Q7OOne2NfyAEx7bQ1KNP155HHY
bDvG5u4hls3Fi9jQA+KkwVfCFdWwEE+FWLVv/U8Qio/9zOy+g6Y8UJhukMpK1Pcn
ao/EDNpOGzuOuQN0UMd3mSBajRPSaeAN+fejBO/39iFq2/SEgf7Hwc6jhdBwqjD1
iBriFNiDeK0oy4O6DJVNfdD5i4qzwCzOSa6pE/3zRUjpVvv2kepMJQrnWXRqnREj
Kx26AJA4LHJX65e3DR8RFaVzGgcuBKxbzyW/zP2EU/GSPwfWUTaPuGWtR0hErpS3
3qtB+EzRwN28ttwoVQonje/Vu6iRMax+thNamK7ZPIx4km/zwO/jNoleS2i5bBzT
w9nRudNMP3u1qZTL+swDWLVPH1MPedSAL09v/O55hWZ3kA9aS1QbGjfaSH6X6ktu
R/we/oslZhPQXIgmkXO0Kf2Q9LYnUVyZY4TWUrlRU0ijMc7UKlvcW1a92+w024Py
ELyn9reKolpsCWaIa2VBAovCuC+QHYWBxZknhxHpwwkngzeVcuQMJgNFNauRgDbp
B8mPkpvlQPEREaccrt0yx2ktSjvz4a2Y/4rtbMK+gBqsXOXk1z94oRN/4ljs8v1H
vamJK4O4/OXmdv7bSGI9Bbu+pEYSTTE20u2+JTOtBQEs8KihsL+Ae7qCxkTg/gQu
MNgzoje6KPwL93KzDH9gb12D/ePLxKYp+G96ipH0iVjkBsYOKtubI9UxbJJJo3KJ
0zHPVA9td6ZLEcsPOvVgsMkI9EUM4dvuJpjyN8sV5GIkWXiycE2DF6GlcGcx100d
FmJdlD9g7hT4194w6731D9iveHFLTwbPvTIdQF/76F0/RDwp8rifptGIMzWLRYRG
uoVxx28pHAAsawey0pX4Wdr0VtNYdmBkavluttYR/vFZzGF3lyqLaWbEJYNOHTTi
LE0/5XBpf9YGgiIYVuRJ7jDl9GNKXYi34Tjdzg84RJS4KYm94ZxmgMNKhWvRi5tt
HyXV44ezzXVialM6sR/DBI1V5EgDXiBgX6Lj2z+/1UUvkTbeu7gvcyuncuHgqbFX
4EkqF5+NaTXgmjjEKc20QN14cnAPz3mQualXuDn5P07egbCHlNQbM53mxV7ERdcG
AaEg5V4A6fxd16FMo2UgvFAy6yZ/tpwRzawOkRd1GMiBqPcvRLDgpRwB+Il6h400
tBgXl3zCKbKqQV/C4K/+3u+Iz4qV7ZAcn2LehBtVrtpPsQS6pyk9Dc4xgi0S8ZiD
Lhdqy+smEArGyc1D8xCLI0vs01akfduKLE4DmOWpahAvadiCtDuJoZg17uOvfaUI
FQk65sne+7tC73Qfhn00Vtt22rSNjcKKnVcvtnWSdB7+W78ZHx6YqNGvyRcAYSaI
yw2KiQ5Z5cUwPzAklQmkN7sIoxOvURufgNyuDX+ZQnk35aXlyyx2dTJwD/KTNKif
pG/uWDpjpUT9oonVKliIDC3QZCI1r9OeJOSiAF6AcTqTcKrK59zL5WQDnQ4qUlsA
d3r72TPk8MSDJCHk+at3K7y3lUaz5oqdkvbJ4sxI2SdPZysFW1potCtYzrSdnVW/
KW2os+76mjYptHsKVwg/9pcW/ms+J/CN93Rir0B97l305hnWhxsX1ZY944JzdKB9
xC7T4a2EokCXiYOOQQZjbUW9V3OtNsPHh8Erue6mW0uduYpHdPB0kgoqeGCZesYE
sHQVAE2P7MzqjMDJJLBIY/e+yYxBxbUvtp0OclPhVVTOAEA9OttW31beWrXDCvfB
OTVBX9jbLZxfc9zUlBZurAVl1YXyJ+G8GD9nKsBcKbo3QEgiyDXyy9PI4UU6qlAW
s2A1RaQ31+EkpyxCDtHeWd7Uo6e1RunMzZskO6ImHtt5ok5TTfHFv0IGMWHrzBG1
ElvZkH+8O82TdOtENsRo3enf4B01Kuf1eTthzTLjG460/KTJls/UsKAkLi9Whxkn
ecQU4PMEVmSFPDzxiB5bUIicsi1qqoDR9H4LmHApRojJ7+lb5WTiE6Gd1w3YkMHe
8JqzKPTr+bcsNfmPpVx7XrjpFpM3D2radQfCWs/Mq7A0Wv+gF/8ZnjumzMNfZTMB
Efbw+JrWmdn0FZVohC5owcON1gMB1tsAn0lkMNfkCnN3kJY3hzw7SfZhGmx3Oz2m
RXycdzS1LU/pU9XVNjnE07jcvZkNSuf6kPZKomrp00HswcxJpGUllvTaDR92oVDv
oFx1TwKOT2z5ct52BVcycjOk6VkYZLc+EYteB4CPTrAjX5bv+yybh1qQ4um3T87C
2qiGW7oZBHFMXx3mUCZAldi5KXXuVHzJJ3oblRZ/NDP6vQPklxU8eUiDQ7dU3mBD
rFFjzAUKXP18bwzGJSV6gyCx/32ubsClAS1wFsKZgHNKPuZLGDcYfSAKB5cPhJ9z
pW7ntWHikYcdxEsRG5me6r+W8stw5A+G9Uw5hFjJmEeBxncGeuTBbdAlujzL/csf
AaxCcy8BzPkDrmrGqI5FsrsQJwuzW1hRrUiY38ad7UvhqbRTU60pugmuR3vVY9od
NniAABlYY2dTIKdkOH5CC1+lxXTEgKJuLOhPpzUUtTrxiVJcFWac/YxZoEqDZfVm
KSXWDgFFzRVHhTmwHwXIE44rC3VqSo5NggV3WYShR1hr0I9Z6xfwu8DJnyTyZiac
NM1JNt9C/Z9wsoLBwJRlN3cGh9ompIYaQoTU2bXdfAn1ZT3Vo4G9nDraNfVPB4b6
mMHo97X3GHQNSzdi3Sp30mpdjhEnF2xyMInGcwcQfgRALplolFJ/qJ1DGhpiO0vM
GAQva4vqllfefJ46FRjtrfkxZ9wmvG8ACwILz0jbLjo+N9JBkfiCKC7BAdnqsK/0
0iiz05kP5TMX5LWxEU3ddMuRILYnjr8DBwL17tREk1HD3CGi6RAPHuSmonnfmkT7
fiy4I+rV4MCBhgk13Poiu/DV17vwrXV71/qqFYqlzZjkjbKhdLmJqevZ0O9BvpDJ
swQvGhdLuu44Un7w0WJSBwCFhe0TPwcRJB3xjyUCViw8lUzkmpwId2aMpsO52K0n
t9fBSpX1IsdULq0EJl2QjS8ouPDEWZQNuZLMRB0jxnBDpcpZmVoW7AgiER7UkmTh
2IQGLGPoLole5PN7tTBqC/St6P5VZVzPsQHCUJa+9IxIWDI0hfEL8eEqtIpixp2e
odH1MFQyacDSx6USucw2BwvyQazhGhz7x7Ws6B2mrFeSh3k9lf3D3drvhYIasMDg
hf3/YZnkcOB5NYo4bG+HvJfipmcVr+dOXCIKw95f5Ks7vMisRU+WQFaxz7u+IVw3
g1NROTlV3vhY3K7uX9Mf4hBZQIx/hbU9LJihaPRuDw88rgIImrUWoWIaWas9flhj
qnimoqSZMWb3yv4zLBjISF7LIogMGlIPa0aoWOWw2CpRUYLc7ubUHp6gycznF0F+
AKzgFfd60mlhrFqJicC5BsrWE3FIL9FQXUWNLpaSrRy2SmZrIIG5+PFJQQWDdACp
xA6Uq+RK1kvXXqohWhiLwBoFgz5XWAj80cwGzXyIe+PozSkqXrajdfxfvK6DDw7k
Pzu5UkH2P8dhw4IdZgJMvLKV7+UWjrlBx0s+H7Gtn+hctc6CfEzLRzmTkC+pvE36
tC9fiHlQskgyYajgODiRwzA2FiJKt585Nxyo0LU/NauuPlfzTL8yH7c8xlxlgbhq
IFyZB2yGFAwd6I41XD+I3dgDOJ2ZIQQHlm8WVIsLG7gep8gwx6TZON/drr/tlaHE
tSoHkZom5OXxDfs+UHPhmEgqly55LdqlyZi5XeJmJef7H6i9lNr3F/RyM2sRPRqD
C+Fh9SXKfr9tzrwnvhXiSQs0RNigtj6YTJ5WAAPqIspZ+ry17wjTsgrUbFbgfCIh
pjCMj1KybvOPRxUXui5LPgtfqE5N14JgnX7QvNSD5kuDckYQL457WWjCDYmQK1nv
/2GHo5WYQrhyxqke7AAfps0PhGQQnoHbBtEwkmYlDgcNfe9BXZc21epSV9LLzG6p
MRWKqKO4qC494uXA0/NgSahIgOFgAg397IaO1/aDgoJ4LuTDongamR+kMvyzh+lp
3FTyYw/w4AZp7JiqiYenRzg/ueI49aFWdHNzDbt9qPh5RgLgA8ny1F4nbWvmujHK
MRKZTIf8bzJdZ/Dwh7CY/rBuS9+Q/WyQTEN06+hRQ5sFLSabuXEPsIORYGhlTkdc
LHo/H97rOuoCE0OsMlTJK6F3X3drnk0fpxdmuP1kup/gY/I31NziINI5gD/t3Ina
9q9CT5zppkrHolqSa1TomAd/aY8NRhVf6JyFoop1neTHs3pZVw+5mU8kyTReqAN/
0xZ8DGmGVph9aaz8zP9nvHhRIUV5mnlCXte0nEOHzFLB3NLlZqa/rHLUUpb0wv/Q
jaDz/gP+fnn97tY9pKaUxZst36KxNct7DA5foNMiEjDQ6vfftWdk1HcYXc+s/dW5
rOnJ3MLtMjCgE1TsGwqbufQE1Bm5QwMo+RsRELkFxAiooEu2AcmxHfEzRgRcH47f
zzfaIN0ZRsVo2pZ4Q9UM4iUG0Fq7TdiyTEwsmKLqZ83g9flSh0ST1OoMsj9qg3pV
1Tklt425KHyDSYsUNJAWg2P7bCrIUomAZJGNdQRshYUy+89MTCT7CVCYLdCbAO9l
qddaenyonuVLnxcQGfk2GxyBFslca7R06drvDwEKOGUoCppKrEB7Waz8qjnLBhRN
pFeKdNn3prg5u/776zzoAs9Fh2cOQj6/HayqymFhTp3ccX2XTzhyvUuYdce6ZiKL
IR1TDEZg9OVKfHSPgG4ZHGRjTFZ1EUjfE5FAvJVS65fUfcqsc7O3Tmgtv7qlQMBo
/X3oud/E6hIl1bYQW2SfLZiMEJaEn9FL4+HZM5sZtB9nM4sPUQO2qeXwMiNmwMyi
Mz/YG84Tcq3a51p6dX9fiyLXbFfo4AD9XgZg3AWhNpPnsRszSaSwAK05girqBNx6
9BMBdi43OkbYqUmKD5x3a5KUUB1vZ8Go3kLsATP/rmfwzdZhmVPHfZ0QCnEB/+hd
IaANFTXsKq7suh/dw6QktNTggE32I5NJvIIzUnOzlgNzIbxAk9dhz5UQH2emqb11
pTcP30NcgSbxb75aVV6z3LJJGxAa12D53u5/Y6wGxnODxwdLUsCvDPpSdYFD8qee
yIWFt9WHfTderawBNmx8YL3zHTxtKV+059kNmscUdQj7BjSWojKqZZakxKbNDkIU
PnhZqEquz/t5NhjHWPAjSCvHEp9ATjLTuDTDUDd9fLbczloZyfvTmA5z+jsofbkf
Ca66bmd1c8ZnVCXv0/uBaLERYIT0gOhnUITMq587algJrTvWPh7aNoPnJjK440Hx
qslosVlBm0vBDgBAp1dtUHTgWUQFLssXcSYqSGuACTxMZ0Tze1bU//+kmK3FsLaT
rTSxAh42/0lX6qjnCSb/J4OAbwv2RrKd+R1kFIv19SMDIiIARH28lz8p8uuNdPS2
blVhHwS3XHT4zRdOVsLCmmyDkWXvOdcCaBdSj2Tt8Aa8KUYlRfbODcpuOd+menLd
tE7CayfXoEnSsskKhBkHfmn7KLtGLjD3YekfHZCADQc2+d5F/V5daY/KGfaq2t1M
yIwttZ25jxk6ON/hmquwBGaeA50R4psiGgIyCV7528RfyBLux0c8iYkS0y3VTwZC
Dg6kLN5NQgoXivFdd1TFSL8Opm//FN5FWBbNZBGz9j6D+pCR7YcBiSQwsPQ2AnA9
k0BdrmvJCRwqVGw2XuF8J0Y+0gtwn/O6yeXHJRKeYXQVzc5UQuMAu5ccJQdhCD9y
r2NEeWxMYZTFGd16t9wGmCCTBCc5DgEEcldJisE+SQsnZ0ed+PVJ1PTJtF3KjCXj
FM8H+FtBjJ6goRCL/MEaFGwmYbNWiNd4dwn404F4OKCv0oKmr0n6NHhB8WjcPJ4h
87g4Nta++sjIJsK+8giWWCb6+heKfOWSnbUr4cWT1m2y0qjJkCWqnelgNZeVO0/s
5XE53qPBdm6rWtQ0Z36gtIFWkMhIqokKIXBRAQISP6xi9ebwwwPhofG2hhmqDAww
Dl8OqeqXKgr9hzwe/8cP8enSe/R6QS6mzRZulFsF86/+DPSKnS4O/EYptOawbIDw
6Itj6xsUGFTYWZit3mWGTodRRXokZIpyvQNSaSGqWm8fV/c20ZWSWEKHrSLQUUUB
CYnyP+imkOyNfLAU08YbQyVkuC6Rgq2zkmUCAhrVZz3K3/O4w+3MvQqdGPlwW99o
BO83UwRKXncuHtoIQrraEoKUQKWvBFqoyz05OqXZ1CeVHNcSJ0q6Coi5A9yH+Rfv
HHT6+m8faG6fs1zmux3h2sebfjwlobwWsJCdomLM3gGbqQ2xCs+j/rnVkFCP6i7m
x4D8p3kaEvvPcKpXmM/PpNFU6NRx17jIsk0vNPxI3c3m1nB2Mqu2YDrLTOxUl7lp
rUnM8HujdcWUYbkwGNE+oQH1FbXGCMrT4VcgxpYRo9eYp0imGApS9M593UlNFAL8
tcFIqxjz7qQne2bt2ljmtzeHii6QLsnEMZLN7Qxd5xPWP6SGQPklfMaYpKq4zGhE
lwCW80fvJFGbX3A38wIwzspXHbTph64YLgq8JAmnOJ47DfvAP1LnNZusAqaXuS1h
uOCkSrDwOqHp8sjrHxXgBqaUqJEJOmJHl98vYkGA0bdW8R2rUsk84n0wd96SI+UB
VbdfbqQ83FaDdXKKC0uipO8EI2hrTgGLU9KSeSQGqPWTYkhYeYeF6qOn8bF+NVSt
Kp1FVWwG4gp3RBbQFMy11orH1iVOJOvrISNEswoKeC8ucyUSq8SyWs7KraJ8D3zh
Cg2i/NmxAkRyyfvwKxtG1rngaVREV8rlcSTM4kC600nZIiz1t2cMqW0LV2PAzvUm
FkEuzRxwH+bf0w8QlN6GKgpjJ9nzBCAxEKqoLUScLXmXPL8PjGSOOZlnH3x1zdN1
e+cDiv05xVFUs4yV84A/nI5IKNBmBm67D6vZgDhwYeJzxOxJ0jt4G1Wr0zzhHuXu
Ibnr7fu3TQ4WF3CccOYl/ewDPon0Obe3oMFB5U4B05+vDCtsUunPVlT80BPKsBM5
pSVmIuKmdMfMoRk9abbpwJPwnTNJL31W5uY48f0qx9JFYJ8L+GSExItqmYvKaCg4
ImJIaibYm2SLmI4L22oUc8rk2OqAPWnN3wcAtnvY4rgxCHXArb0wmAQxB6Y0kpxG
WU22d6icF9osOwME+19wx3smnZuE+5tiV5py7YWjS6+6r4x9gnotHYh+Xp3GdaQk
oLJUAtKFdpdb0J2tpK5O0Z6Qv2wWEcRleyiC0si75qpMp2Rfs6NtLjOvPO1lp2al
Be3P5m2wOvFK5iydXgdvLQeCu7q/9FeFkvRAF7CNVtcJ5L+8rO+bLZt5zf0/GMb+
alcVl8WhfbGXSkpG9g8aQJo8QgAqzFWYg8WJAKH89+mNY168BV0nCbGVsvDeP4LB
zVlhhYIQhqcu3Mkrnj/xI2JMH7oJapx7XATES+NQgMqN3PWEOMy+VLjeU1WoBniw
U0Fj1wt65NNVPTxvbFtBh/VGGiWSTlAsd2OXcOQ96tTGubwFypXm8JDqhb6Htt8t
S/TDziKw0s8xb4uHtCTnnEPuBN9qAZVWpb3LlewiCcJe3d31heIvrb8sxCcrBTdx
8CB9ghNhQpOPvTfaarR4608nJq7xbVZrRB2uNFKDIDReOpLMarw619PmVnUMorBR
idBt8v9ydd70ocFMSMT8rNmvA5pUVfogT55MZovZshmRGE6I35AJhJinHUpwVcoI
iI7aRb2Wm/X2F85W/v6h2mnBX7a/ptmWLitLg8tWmS7JphAOakYAoT8DhZBi88Ai
9+DsOFG17DYmMn+n7yhGacrjgFMGwhUsnpfJTnqnLB1RBas5sgKDr3cJ4vSbNwP4
Ml/f70fL6KtebpH8UXuX0IYnAmSlZ6xZHQogbVwBeI16BNg5kQfgQAHgl/27Z0J3
28s6rr9ZJv3WpiL1FE1cnma7BrDe9hdX5Fw6YAZpWUNjv18BMV2dluS2WkK7ytpx
Iv9egFZ7TeZItaq8U/2Cvvy2EE1aTfo7Tbb+13P1rM8tFUPcms0bvd59tik1kRah
sUGWuNdTfYZGTPldHFPRtZ5r6c9hXaFeUmQrvoMXPkrhtmO9SZfQ6wiUMfmhlsBb
VTGDtQYurL26KkB4KLeoNerzhQkVBLOOGVLcTbEbx6z8fdt2fa2DWUX3jzQ4A3SQ
2OhwdQJFBRol3UAAmlaUQqh8dRfVax+d07hQyaBjQmvamAZlhcabVsrba8CMueN6
B7A0E6DydntViCMMCPs1as7oejWvG7U2SCh8/AhW2zc4DAAMcDWwh0tpaw7zSaxb
V4YBF+ZVXzj3I5CRkBzI39hwVGEaIC84Ne00P6mgRvlUesLVykgXzltLxeZ6Xl30
`protect END_PROTECTED
