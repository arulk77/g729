`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJfxZBYFbXh2OoWvInimnrz6EcAwzF/LiTqJCg9DlPjr
vsg0wzVK5mQHhjbhMNEwyyqf9tzJEs9HNWfrp8gcMJKyMkm/kAlAHntxyJmETd8Q
5ruxNLCRtC3ry29mGmCn/5/6TNlZkloXjK5o2imgigHn8Cit0BVypeKjHrXZuX1v
ORga2OC7WL7fvxfFSDXg1KxdR/oXno73meEe3FPIot/SF93vDCIJ0BFkpE/duAYw
1q+zaUOt2atVNeJyJuJUaFmfUMK4ZXjvJxm8PwFL0JJqUhF+mqUPkgOLucttDt1/
4WYuuOcLKH0dgIOk0s1QxjtD+i/eYMzKNTuoo6f1QWzjU2EPsf1R+Io/a9tM6L/n
`protect END_PROTECTED
