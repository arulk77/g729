`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDuF0gMs7IuYFc1YzoOkeUNTx+JkW+EncC9wAoo7GD2c
y3Q7rxtt6MT3ZitA7/OKTtsKqlMD6LpG8Ord0VLVvkWA2BnMrDMn1fawY5gkKhD4
+clPG9doDZCPFhNYf4oTfcyoREhniUEirvikPYAU4ku5+q8n3SMldYIDu+vQYbup
SODxypdfvOr2EfQR8M/qp7Ulv5VPDKbKXPZDGOjnwdOOOjkOoLiuLbdWezOPbLMh
pmfQCtb/kB0DffmhJTkKBSXoeuZ9+PFSHjnVZ/hJmpp85cSDPkpq4KpStMZvo1B5
V3gcveeO9l/zRVRnZwzXmxoLDwgMIHhLOb7U6wfr2MqdUNi3nv1npqW/Oethd+hj
GxFeNb8/T7YqjSR+DDhYralnoVLAApSDJyl0449wql5vwG4pjSlq0Lh1NR6pOTGD
AJ8korirfowcSeVfQF7MjaB0QQWtNg6E3RyXrb+YYnmMlSvE8lQ29nja20cRYAPq
nIdS1lXxVy26emOH5cpK+NOMhh/zAXaumLoyhFD5gp6khKS8/x9uwn8o6802Snju
QYSsrGVfYQ0GkLNLJJRNUO0NTkAgf3UYpvkT2QGQ/MdeeyYvPJvygVk8SFUPs/m3
XnecFBvVhdpDFFnOHv6nDVPudrupg7CWoPnAJSu+tcs1jEz89mPy9sxcHudfEz7+
B2SNOV0IVBgzhR9GzuFMxXWtN4y3pSp3Ayk8bKySEk55V+hkg3vl2Dw4GFnFB2Kz
QagtKiQgxIaQ9ZGDry+WCDEeG9D/OrO/UXeC+uK1kkhHeEhXuqlOKszuPqIhhYIw
9dLwF8Yb3gef+kHklHg51VBUlyqZb6MLD+LbVjz3NtjU5ElecWuTxRnaSnasDpnJ
P5kK9wnid6g4ogpW0mBv0HJ/pFpPRJIs5YoygaUp8ZpzP4X6HbHBtplAoStbFK9t
`protect END_PROTECTED
