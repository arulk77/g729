`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NiX54RfypJ+3XEMWewlaN+mKq5i5wlNKNui5qgJpZ2ren/u5ZYiiUUYzhKgF4uMo
9NxN6gMBtCeaAA+lnJuTC12kCynrqEkQh9PdDQ8wSOX35C3ud6C65r2Be4zEwIRw
qu2I6gfoA9QPZAFfWD1fQZ+X1WVwKVF3qU7OsV/lF+fz7I2XisqiB6JVd5NBmV+t
6zn6G4k3Ndo2YADRyCRxWbpjEDLsZqO/8UogjlY9ffgdMlvzSsYXQbSIUDDgkSDH
Iq4auhKCDCQAMJKPdlHSMJjWq9gf3sCNVYVB1JvYbr4gtR7KBCN42OiUc/rl5yqB
29LtCaFxLhDXDzGBeYVhrQrAXYJvjlGAb/6iWrN0I4n2zpSG9/NHXqC4iAP/Fu7m
Uj1mDhlZPHQdB0RPJYhuDSM4ZWjQRG2wUy5hMga8N3GT35GL0S+2NGbsiSgI+qPR
1xeKk8cLk0JE1N3YytEJbEFl48kGnZgpNBX7G23mcnI=
`protect END_PROTECTED
