`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46NpC71W3kX0fkgJz+rEHfl5eX/FDU/HaOBAHETDKSXf
99HEklqstN/cwwmGAY0awnPpPqY4/6jwajaKj3rY+TjKISvn4xB7atIBFVQsNYt3
7bQP0ni5Wq2KI0GXiFonl1WDnVppucdW2UJYqAgFSWvgHMts1f1OmFkONq7S4YSB
8DrqgJU8nP35smommBmy6Il9Nl5PADCD2LmkSKeur5X8/pL3fBgA6U8VkCQfhofB
LL102Zdy/OdsFnARYu7BKdBpmrWeECvh3e6tDsJkMmBdnTTfQ4Dc+qu2ruTMfocQ
NgrQNozbRVRU1WKmhcZPDQ==
`protect END_PROTECTED
