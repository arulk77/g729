`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CyZTYWZj0nq8lkyqCcyi22oSD5uz9EvvsKWLrDDKfKBK
6kNyTd/M0ydoKX3W7k4d1yByDhcTxPEzIZ8ZqtOCdYp7IGJa6mr0jMw1Tiw9NsrQ
67I+O5R99chGzwVLm08u4FjI5hDFqCkxdLIK2dHbSprT+WjtUi89NfYph9lfj+ol
ckJs4/bWse8eDWOBlt8ShaLo2/IlwtdheXpsFPvQyQmhqEQ9FDXf3kREy/+alGcU
T7VzwD+4aaDnLy/2h1N0dIBKTa9K/KjiIaC/H9YVNy8lbUDpeZtx6JUBDHHWq5F3
4tvDb9UvHYTjnD1AlXq4hSqwmLv/GE5S/N5qPD+4ZbFckjR7gHfOuOgbMSNMgUga
fiqsxcX43UoDG/JEAG2SUD1hVdGbTkDeW4wEe3UqRWedJ9JRFjVu2njJG+MVnKMQ
GB1N7Igij3FpmchkVYAk/nr5tPtz/emG6AqOZ+spn2w/HtfpqJJf0SSkoRm+ZpDx
AK69ndQ/9pT1dE8Yrxy5gS/v7w/eSxM1TEzfOWydbCCjBC9CuEhXcrDcFwNIQh3k
xnpQNoS56Jo88G0nxoNfsuPTryyd/3awa3Iv40NJV4J5gkwijrzXZbIIC+/fUbQY
FkSoNU7k0LpQDHylOk3q9s4EdXnIPplzncSa3mb32RVE7eb6HgIK+SFRXpvfHwtL
VwCTDhgBDt+ZKC0akjUo2pH3cKjQ1OMvAaslZF5X4ODarHBn+zv+ipfGF72c+5Q+
BcUTOf/vgFFFuXJuqlA0GowS/fUNVp1WJZcZ/DcxtHH3zMmjferdu3k5uHAC983I
myIcVI7/jhHqOa7E9gwHwIkvQ0PRJFc3Wu916Gy1gfp16DAPi/Cn7/UbRwoYU/eW
tr/h2ocQh/InKDmByM6GVi/MerTpt97NMjZjGiBe7Daib+tf9r+tCbXV6mzuuHET
nFXctglQv7TOjHXa3NWMO88Yw/n3hZ57UDUbGkFfGqcE5vdFJxcjm/RokYqYBfOL
o2A/hdGp8yKF1LasUMoTLfUQOvPZ9ayYchY4v5YmTz3jcsA2AnsbHVAWnxFBvCYr
ac83wSDXG2sOLXBCcwkkcV1xGajxRQncKGRX2vcr1c67iLY3/IrxrmFJzM5LZ7gQ
gF0gzeKicgSBgkiy1BdJFGn9OMDGsb++ZmdmCHQrI20MuDTPEQqxAse0h5AirX7B
kg7CpEmdrizJIIYGi8A9NuLGW8dvuiMnFpSJF6UqFGJzJdp+BeJFx8I0CF4FpdGW
Jbco5OFKC8R7ioxTRR4eee3FwIdg6PzYah12x8J6ttRZ8hzPbASXM+PGQOaJBjVP
w8GZM4LRaKW4mDu1PtWJ+Q==
`protect END_PROTECTED
