`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKT3CMp83Ejtehkm4jdAj/bCILMEQH+RA5Edpq6qJUl0
q/uwCXDXNvgE4UsI6allNX4XGz8ufmjyLWS3T+nBIT4vWeqo4MIh5LXZIi9VTEj0
9jUAhRW2rjGiNmk8umCLRcjA3U2snpJrvZ6lXBRM6AxS2+SBb51eP+K0FfRVIbWJ
`protect END_PROTECTED
