`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCWSyHQPefsbfR8U0gppbRTU4zBbwf+o3xphYrdJ4nnj
LpLnE/EOBxxDlkDJlEAriPIdlhwBKVG+AkIFRvvOtH0uV4KOdKlEbDRoTu79d+r1
lL6U+vSOlob74/HSUXBC5M602u6cxEpq2sJTrMaKJRU1iUH3T8iharkvjO3Rig3h
90vUjuiuvZcewDbXVIbPGDn8tC9a7ycb7pJldfu6VsP1XPFSy0SA67Lp8QAldCi9
BEBacT5hQ9oRaKtyY09QsEWw0/MH4U6WINTbdeYzLmLYcWMo9D8d0Rvf1cz1Vnms
PBTUFgNBkCMgW/wrolHtsBum1uU+k20S5hm3sq9l5DUr9CfeyQWRh/q16Npn3dIz
2VvkKcyg6QcUWESOeEOXbmELLsHNecXePtwrmPyRPVNEBBd4DjH5J/a+JJDKsmwd
`protect END_PROTECTED
