`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
z8zz5Tho1e5b5oJ9Ksn34LVmvLWR1PKSG/BG6dQZ4bTdzyocHGJhpVQe3VZWRkGq
9fPWDHesQ7zimNI8QiF3Z5RPGHz7ZssgDNXmVFa6Yl97gjWKepRXJneXqwcQIokV
lWT9QvchlJG4UBzK2jLFunyWyYezMSJ+TxNdT/OZyeuILqoaRVaQ59CKcfvCzjdy
`protect END_PROTECTED
