`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBx8MIizcw8emPdE0gJGSZLRYUw+Qri/JLk8Nspy/RLS
1YvW09S87e6TbeM/ZCxAmcqkoO0osw+MARTv14Fkzun6vFy5xPa48d5DihnYvkDL
seelnOSquZlzZq4sdY2SPLATax6cZpAirSsNCNHdrfWlUjJpWYRXeyDApdWONlt1
TQMp88Co6wLtwEtPkSxzTTavqq5UoxQa57IL9lPdZZRyeI82y30NK2Xtj3HDijbW
fjtZmQp/zIMBM2yyMfwhy4Vv5HyyR92H2dhxuhJ34FvuZS2WW0t9idbrIvfC8hzN
ys4NlT61Tm88RVtk4H7Z8mTpna+Oq7KPNS7zKJ3sG1EicO4wfZO94WnwpTb+8Q1q
5oYEj67n3AkD4V4s8MyYERzJHiITU2lnA45tjRzzIBsOYx1oRYEOEna6LRABphXA
gzzbUPTYhjSk/qTPIPrGdAqdq98mqyvkp46YbV3AFdhoeQlMLUzES7rvDsD+Uz0k
Pp7SpJyzbxiDZz4ZLhaqy/XjLc9SKFAIZLzbjrVtaBmjXZYPA+QeHsiKWxL9RJxj
`protect END_PROTECTED
