`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCzpC39y/yxIipzo9sMF4FdGe02a4iZ/bKp7zreSeXUx
G0NJdwY49ktwdtp2rihkkt/92emnRut7dTcECrbtfPMQzEu0D+v8gs5vAIw6Zlad
3DJIm1dm3q2xU2iDgVBatvy3SqvvA0lXL5LL48TMk02IN7PJito1Cwr8tuNKx/Et
zqLVqBRVEU4pTx02sMa6oshPDp8O1o4BNZl7C1OjC1/x1qhXA5fAZrXZRknZ5Ojd
5EV5QvpJ+hmJYxVWZd4q+03q+W9U5w+G0Kecx/I4lUoctqAGDp0DbczOO96fYKog
BzfIEHxsf5yHLMehSokwxg==
`protect END_PROTECTED
