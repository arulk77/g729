`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SWw+Zi0Iuy1Y+uQmWrNeGFGLG74F95kri3H73C8oraPT
L7AZQWXX5d3PuduPpVKNL43QW59hDZBoYA0NWGC9aWxluGVLxYQaB/CHxMyIO3C7
YqCIKthegs7EaGE6SZIotbkJS+9AGnMlJ2D7ZShrqqRb+ngTaxvZdEAue4zdnlnI
qKXGvpsfRmJPy7uarba6cNvvLEdMrL3LejWmv7QNy5TU1+Rt+ZvpwM+kgf5sg/KT
YAuasZEwKVZEOfqqvWPN6wYbONVA6FFLgoDG4fYQK6NpvIr+Mm1aQSHULjBRlFYh
TqggMHlWq/e5Lw8eL3UetvPHAhIfeDg0rB20f700VcXGnXLGbl9RJut+ilxB3j20
n8K8BP8wc4nS2tDbzWXeHXOopBi3UAT+FNglCrItY33Fnvqq1FK+10b8vK8calH5
TswbxHq2tRnxqA7aZ8+tEL7+HN3WfOKjQvH/0BWa+1jg7DwwKHOx76zJ3EMHCbQ3
4yl0xu93cQUweq6p+ykBzA==
`protect END_PROTECTED
