`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aV2WYNgm7yptsHIp2C6YwdTfTNcO3qULEU4/OTDJXIN7
8bkL4bYh9a5Md524fpNuHImTlB0LP3tohmrJ9vp11zKaVvUi/EJDnKD5DcpUdfjX
eiIL0Fc7+RkctWVFZvvlW0dJeAh02XXgtMPt/bWaciqUWI6k55TXtU2kMdGIAkTm
T2GuDgS/mZ7uwOuzuhDJ23Mw45wRVd+bOmPcPPW23H7Xhf2fyFt+tiWC74pIuCbh
k8lF0YSaq4ZFNnJJ6JFDCFyqvU2yeeZrlPXZojk625yDoBhEUu40/riV4elZDF6O
vExirfy0dTHh//Ec8SXP8Fn1XpraPeYLKK5T13fcvdzyJRm8BqkKxt26mPm/9OAF
AAEAKQ34Awwa7gIqpb8Z7QYkh3hgN/qtQTc3vSVTc2mjF4YWMslWgYC3nb/QEtRO
7u8CmU71/M6wxvgf4KeNAeXpduACdelr+meQ6xBnfFXosVQiz+Qh1ptNRaG/069X
ouUL1LY38AmfRu/Pbt4faEDzC7O0WMDPLW4slGBGzLPBKwr2DPDrfHexlDbDJYe1
p+ldMCOJyfqBLL+IQRSeoCUVKXCBXvsOP+hfhF6KQ6OZzt00Sm1NKx+85v1csveY
RRXry04trpbnSV4FJarTWNrojsQ2XIxCqzeK/8F7FocTVfJR8mZ3CvhmLK4Ih+U8
ziYhE1VF48ufBKFAHB4ZsQUmALkl3rjV9WF4QVjwnJDbgqvYLTexkJFg+ebFE6bl
iKn0PfJCmaPXtFHAQiOovoTKRM0UkkVwqaOPfqanyw8r/ypkRT/sUlWBFUUTUF2E
xaDOsFIW4p/gTQhy8P0kiCKT+PSxuhZHHYDERQU5+dQo+VHZO44oCgfxcm4fVsZ7
HPNJ3f8H8WcDMe7m+H1hz1LNloRBTn0QIZ3q1GktqDAZKigY0uRGOPRtNzWCozpF
u5so4ygYGoVPrRy7kLLcERwWuimU+hNQhk5+Q/EHYxbWBvNgXDaBOd9n9IbN2Y/2
gudYwY8Ma8/BLANzUgX0e27mEFIe8EeBR1abUIU70LasOwY6VH05puh/JbQcOrxw
fKJ4Co9Gm85IHvj1y6eZkiDhaQ8N+YjhrSMZFQm9MEFzq8HVAh2UDKM+oBiqUjLX
vgKjXQwKBlnrr0avqtXNUHxgJ0ivfTYkrlS5Bf57xpQsS/eXe1qXOorQh+a/wP7S
sIME4bltYXy+BP+gMM2j+kEyqMWCNxx0RQ665qLwIwB26Lt6gY7pHF+dn1OQq53Q
4bbM7FNQv0tdg2fMUzyMzo5JJQLV9J100PoUHi+Kto1SdiVkhr3jjKu8pnLEFaEy
MUJiMBbpUXRFEiTObFNikRrAebizEILV5wTdeJkeqm9RdEtApeCzZMg92UEXpHGf
h3+8QeECbRRS/Jb8bgIBr31mW1gIZzYcpIaILgTMpc64Z8GzEi46Fi8RdPfeFgDa
iNHAWSAZnTixZwEfBVjOjoUMP8zJhlR4MemjtyuT37s9vQ3OoD/DvN7RvdH66Qkg
yvxmrBz10sikDB4UC3KPXIp+PPftxOMeodkDOFsFpG/iUzcljw4HorOaLSiWjihv
268itXp1bCgKvrRLky5rbbzagOByIi46r2dk5NjExSvotpGbB5rbA+HmEKns07Td
zX1hJcCsnn7E28LurP5NlTG7SY5IPaYuGv42teUnx43hNoCqtfKk7DYdATz72hJV
aBrVdEiAhDlHZDpNi+8m5aNzf09/ZGj7QUTVFhav5Wio5SUzqTN8ShcsgcIa8z9t
1c6N28gdFxLVxriHrNU405/NMwKEXmo3CpBmvd8wnRD/1bc43HaiAh+2ZhJktrDz
zFNdSXhmhcJFloPrKSiC5S3PH4L14f3dW0EazdfcSufQdNwmYKKc9SR9Z2oSlAhd
W9PPPwYCIKG07eChe2Yxx40DzB6JWJ9FX0Q+cBoYI3dBx/njYDAev38fqy79v2fD
Rt+Hne0gigVww8D2d7DfJ+oERNBnH5EekvPxVGiMpOD1/gHJF79J//Ge5MoHmWco
coI+a870N76lYzuISB/KszilQQpwtXKbcXgvJfC+Wmc6aF2jiTnLrdTc2muBurzU
YSK+vLIa5s0k9P1FQq0nBWZ2RBQ8A6W09aGlxT8RsUuie9Xt4JTh7YkEblfnQwC9
MaQpuFiWjyvBhwbD+kDd8oqp5isvos+5GT80195vkKSZjZROXuUTvMnLVkTx5e0Q
NJHauRYtS6/8VUwuibBC+WvXfPaOYcDDygh/7IpAMdgKlEa+A7mWvZKqjUS5gvTG
F5Htoao6XWVNEkYmZFI4CYWmq342fxmDNoi8xhMwPfoNR9H7pfFdApRj58r/yktJ
0oaIYaOCAbxTSYCGoek7VKlPi/sdDzyPBj5KvP7KV28OtC81IF9rO8pRiqOkV4+r
fJzdczjLL0i1in230RSvMwaOjQJj+3ql8bG7BujvBd5jF9UH66f07Rnxzr+XWpcz
v/pC0RDZ4Ps78kncvMYp/gvIdI+3QKxs503C0LUk2XjtkxJXOLxxRvKltynjirew
sxRg+Uj5YslMdtKLphv3lZHYejN+uDl7nvpZRWZhP/2ZrAilaOEaQBAsFZeRe6BV
FE96RISiqJmCnAdl04R4yEevfW7cpoZ7gbkRaegsqwrFeQqgq3FjKZiiXu5cEeSU
NniZvRtiBT6W+QE8gOn6f7r3BdT44OuvY393pAwoIqqJp8S5h/Ftln6khobjJZzY
Aahr+Yvpa5zj4CFEa5J/kXOVXtlq5mVhfFvFKR2L5PiUgBldDlAZcWtpGgfHeAiN
xDeqUWDfN+AEUiJ9Hacf8KBcTlCANx+Rt/+SwleagC16Zy9uMiA4YCfpxWhInsbQ
Iui9f1em1YP+Ub3NH09ORHviZm1cmGBWvWRS3r+XRc/ILvBNd5yNqxTeESL3uhv0
kouUeOuwpoKs8sDfoVMp8ZxtUb/4mPJ6X8NdUaBW9UJw7W2z6tfCm82RLfLBzScV
dOOevKlCQelYD00JmPiHrO8KWTlM3WN38iMht20Lfz3r/poVLQCXYCqeJEbetV06
BgWjIxHEcvmKBDM/vswoAZ9CS1UFN3CsXn8/W6wGvnVAc/DhRnffmWF7q2nsfsXA
fn2VRDvTkWwV9WUc9BAvWA==
`protect END_PROTECTED
