`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEqdzDcHPU4xB2L9oIyCkl9DKEr6sz9Mo08UcAFRQ44z
o8fL8Rk6o4OODTO5746Df8DU+piGIphyM4kWySQj/kmgacZqO/T91nRL2RKQg68Y
I1AgVd4tADmQ0bOrZZkKXBgOZNuEPQIm8gISdB0sEL77dLvG/AuBypQedwB/SMlr
u3kPGbZyZ+NXzkRZqMgZBquLfLDlt+NHKPdYdql7011XxdDkmZQjnwG48peYD213
VwuCsah5PJAaa35Xq+SAPXflK8Fs6EDwwTK1vZ2m5AZ6UMu/7su7YQYBYcXTkVkx
S0kkqyiWFECXIQtATIw3HAPK82WBNOEKPtcMC01Xe7NoybMK+n8nHc3if4vTJGOk
JzG51w2ZxrerYvyno86JLQ==
`protect END_PROTECTED
