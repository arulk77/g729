`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBM/4R72vTvtQsXI8HogORe99wzpFFMGry7udNmAxFXm
btRwZrYE/jkjYN80erSbSm3qgve6kxOqRReqEQHXMGvBNhc1tcjGy9QaP0xezavR
rreZGsmZbK0KEP0uF5oUEPg6MCcxG6QIoPH/AONrduzE8tUtrST6EWizELbFhN9q
PPohSzh+dcKY6FzS5/rttTkKLCtwZRmxeX6c2kc3u2yC31C/d4yZlLJKuOP/bemI
1mnCuUq1HRHgzAVTNy33ipVmB2cyTpgh4LhyQN10uXdu4d9/YHdO99XuSGZG4UHo
DOlAp4k31tSWeq1stqhBZxttSUFWj5fIU0O1wVOIW1c57IAMJ/FttHSLD6AjlcDQ
7P2TxaoC4yJmQNQblnBb1zaJp9FEDaUGOn8G+56owWYjQ0BckxskhcKHUbLbLrjj
aKYvVYKvLvZCWB1Tz15MAIdOTU4rEM07rUhr1H+cFkJ6Z/M2QDuwkZ/KZJfcOmeS
PXKJzISflQ1LAomS7yxVB9gHbIvrguaPZA6qB0B4ECgylZYKM+aO+eJRTzfgCpUf
F4ZzI2llywHUtwxv5wxMfmdcBigU/mm/RbnuFEDmnXJdscORgdcYQNuSEW1EDek7
Uxfarlokc2WiusFBpPnT5t3KR3eqLRsRubcPud20xCeOkDqXrkYhrWvpN3A0VDVn
SpDYEmK9EQFeNHDnwSNXijqksjH6SgSjRZbNfQeDlTB5XgR1CXx6H8tpe3yVCtj+
vJKp6mxj+/2ZO87T38hbZIyf2N/y2HY8JCPNLKNmtl1CmX46pEBeNqVvLcF66fXc
RVsGM6O6IFiw3/3zCLIT/CZbNyTHc4CADlMtxYHAwBW25a6/scI9yyYgfA36ksCF
cA5X7O6qJRyw9jXUVnz/3s/ovSTPGlScZ+75TCFU4NKtGHaVBqZn8usEvmvCBrhH
h07sjWyPNsoUwRKJhTNh4vQ8LA49pF/RTodWZjudUlp81EVA88BMiuQJqZcisppO
/0n3K5NspTDLN32l0jabtHe99Z7OdoxgcG0MkpiSr1jKZeBXswXVmHjvo7pc8EMC
U6HYTKI4KZ0FzKOrCC797O7AAI/e+zH+QFrkv9B21t8=
`protect END_PROTECTED
