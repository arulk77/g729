`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZscjPHZzwrApp2lUrB0P7a/8mZJ8EBsht18dcXjs4KMZI15hhyM5N1Mugr0rVWoG
NXFf7xyTO0oBIrPdZPs1G+pg3aZBD5zqT1dIwmvfgE+0rHDt8rY8Bfbp/M+auJ5T
14HrkJrFKP7sW7MMQDilnwjIvLiDLbdv3urHyg5bCeVq32IlHA6xmvpXU70gLk+V
5fLCvxJ2lxvyMY2UC5Lh69741tsIhY7OvNrQ4/4M3k/RyzOfPOvp1/zmEEvgDs3H
kg1SxA/5fkQ4EQfldINiGXMAtEXA3F4T81tFrVXwD8Xa/KEMlzSqt5u0VafKrsN5
/QkgwjIYs/NniEfu54TvFkRa4vnXb2+FMdJ5dcLRpkGjVwy+8UMdW05GEtFE3CL7
jIdIjY8xiz99lq/0dW0yGb67O0mbELluvKQTeNzyADb0oVxO6VGYgjROXMQX68/h
Vh0+gvaNL0yvrihYdKHiU/efHROsQuewZJZxs17tRANzozjyX97ufIX0a8uPmC4P
MYHuk4IqqpiHApVEkq1HLcyFOkGWMLIi49L53SSz3CyBgX5o8l6uHPAJI92tiWgF
iNaluTnwoKIRthICQ/1Hd8rONWDW4tt8yqiZAsO6KxlMwqowDXlfQBQH+6TBq4Pe
4PxykOSmYXy9Cc0AYuV1i62RnaurzwQXChUiGKa2HzYozuOE6sm6x/JAvQ1aSw5T
2HFcoAZsrZ4cSUdOKuSgFzkCm42podjaC0djlguCc9UvhI8jxSx9XY0EFaUzlaNt
joJ1hav4BvWgAgoVh9kII+YdJRB2eudYIb6de8vfCaI=
`protect END_PROTECTED
