`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD2cPPRZnVBJE3SbSUPH04YDBgXSvKP8nYQKJrpENmoX
C+ALQGvHLte/it3x2EvtbZYB0bAi0koC8p/zuh40mvAMDWheTFu3ocXHPJUjxS2m
4dQPEJXT9DpyhEqUeI43dZ2t1GMZQRU/IdqdrD7Le9wZgCZ7x7viGlD/aou1x+ZY
Tq6Z5QybID4ftimH0qw+1aFtsj4PjumYTujibdR+pQQ5D20upb5ccdHoyIMPbFyN
rsHuwSiUCo6RHFjI6cI7oE+0u4J2/xc2OsrJSThpOYIBPdOUQgIb0DPtkKKMpkr8
tdosNhZAX1OvPdn8hqJxaoYFwQyhA5WpwA7VB4pEFl/GEqIv83H1RcoHzRs2r8Se
l3ZuOgQIy+N5md3QqG/zS4fzrpFlXXxtYW2VJS9lpTiH821LIMWJXCBGQwnKfatz
/S0xmvlJcYSWB/nnBvv8i1dnJazSDbK8A65/UOa5iL2OcTtcJoa36YAu1d/1azvd
O85BAZCui+ieT7lowavI2YA4HgTzhjKf272rLD5BQf7gJicG36qTjuFhbB/2gbJ0
iEH6L8hpliz8ISYkfxsJ0CzTYOLNkKYdzRBWaTe+++8nlX/XEwYN4d+B9h4ibFns
FLUVei73g2tBevTIlSbbHK4khdhLmgR24+qliFBqw30oiLAUHmHVMfBDd7XDy3G9
U8Wry4hxc8V1JT+C85kTOg==
`protect END_PROTECTED
