`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN28x5ncLRDzrsrx9h6/rd+QRuyQlRyJc/XiSFnKPl6xD
QdGD2n4zVJyEi0BWNdfMeCYfkYjeCQMrvY4e96g6WmiHgQW9pmMoO0aA/WlgRrYR
28A/dlfja8zEdApf5GVcj0FtyyVHZuVD5LOY/s7P/BiKOH8uEKZJFi0l++qcrStY
8W08PTjcrAaLcCvn+c+dIBkgtm5UAF6Roc7VlqeheBONAI+kPCgIPorz8EaGC77Q
ohqKTXOpp1rbl1umrozWrl5O9hX+XFWOpcrcGJElm252qQUTEd8Yzicu26NePAxB
aapUXUZHe6tpnSRmLTGLqahYw6lKnfye5GuW1gmjdpDuh4R6DwJrs2T3AVW7qhY2
TqomSoEeswG88ff/aLGKF6VttW7Q3IImlnciJNHqShxxRvTzk2qRHrWJXZB+fKXm
eDnyECRWCd/v+Ug8QLf2g0RaR/iPUO6lQmpzgYLVlzjO7BkLg/8NaMfQ53dSYzBt
FiVQF5qSP4MkX/Bd2Z9ZG1yKbqHtWv8+cYrX8yGJs8MxBak9Ct/j3jxMTzkMyz/V
3jgDY87rH6jinxBEfk5YBTqJ+M+2pwwIGt7b+3eQI0un5LhbJvKu+VMRScAqRaan
wca0dqn/aw3w9/gvUxf0ON+Ut5pgEVOh625xy40zUob5lOklXG23hV78jHj70kXt
N/DRTn8wlObDoWwjZrpFVsHo+pDN+7VRLsFYzbA4aYwSUeF6o0c25ZoJC5fo/7VR
phX0uFkZ3dYI3IUNNGsZVzMvRg1bwGdJ68bF7RPQb2K7AYm6DrsJCCmXhf4/MMLG
bY4tK65cYM4hG8BT+PScwFN352Oozg0xuivrlXkZv9JtQnRe8FXWVSn8Oly/GcSX
gKWFvl8tFrGLkqimD1/JK49DgTEZ7ndrRfRS8enjrYPXfSAwiE6Y5tX5IEtTqAU9
awgpeNSoYJEnT7jteUA2gv91PEwHDfiRCeAl36qatMbLoG5bF4iwczKhGNe8Tn2G
vMlHbdc7ETOD/PmBaIA1N5D10armezZATnaTQ7AWxqtVuP9ZS0vJpC5FRj9i+3dm
aZVZk8BBKS5mriqBddiFZx/uX2nNNx1TgoF13xf9Ilr5nbdbQDaHD/vzdL2+tZ8G
IOq/jqVCslvzvUUuZyf8wC1bAh/wCUx4XsECaC5P3PlELdlp3UdeYZDd+LXbfAYb
NHE2I5z9u3s0C3HW/HMtfZc6z0NTSWJgEhoiPTxcMPEePsGQa0w1lex/1S+3eyAi
agD01reX5rfao++UCNfhJByB1lrZRdWnLYiOfNDGMShvE7HvpcopM5lcDyoSlSih
3w5PnVAvg7KV9gIYZllyopI9ipsBzjQ0VGtFOWrPTkEKjxJOj8IVrfk5S0bDx2Uc
Sr0YOrBbcgdKcCrRFNVso0EMugUW5PwQCEwSypDfbvIhEPPuvhxuQYPiyAdtZZGE
D0fo+hAmqgiz2XoRN3eMyS1UY4JE4PGAWIZxHcvn15ZxeDMBN0evDYxNCSWBqLi6
nutzz8gXKbV5ylkHy4D+PPZitc4cjTkgZkrBTdxDeVI2kgf4+edcXW2/rlFR00Q0
HZvlcTFk9+6fOwkBoVD49A1u2NHZQPwnsDsRfLuaU056r4wr7bPRCjtosk/IiaxK
LiwVaBuQtaPgs4plzat5BxB9Q6GYsrN0KPajcTuI4u4S/iSBHMsxlIVQTbnM5AdA
BQaBDH9Ao8u5O6F3NvyT1jD7ZJ6JAvTnmOPc3eVgXAJ/PV8/EZr8G9bUfcgqZ2aN
wfEs5eyvk8KIcKYUTjKwREGo8SEjLamnaXEa4SRPyrjSWvxvnsAbfDNHJlJKLUsS
WLCPjHIz/Lzk7uoI3pUFt0iVBCUa1RNcrYcYtVOoVeMdq86FL0fz40p3O+T7WgPp
aZXaAe0yDe9ayS8Yg6rsm+JQNdYBiax2Mum4EHDjdQiopZiONjXuOQqFKizfF5Xn
HU3hSWq8qE/+k6vaeRx8Wx8uhyQUvKxtma9lhk7huHrD8m79KWpAWE5Jo8f8VTtt
a1fqNxhE5YzD4G4ITlhXQ1YOrJWgYbjXkPNT00opbIuNapvzdjCheqZO9YN/k0FW
0BVrmdmDlul/3QV7AtA7nzb3jQLsT50L887PfkUexHJObUU5gPrHg/S/VwY2VYno
OcDFlX4TR/svR8D9XXW9s8R4BkznuTN9jg4N/bi4PzRXhYhve1/UeWXuGK+NrLXr
uUtgz4mUg3flN4cFVPAUQUxKApUTODps4Ri+EJc4+bGDPKX6RpQH73qkO0rnN/uE
cwrrR0t0S1qCDL7Zy70nYQ0m6/AJDoM+MGdQVlCaUIaobO4TxDkEqkNbXnwRH3rR
Y4NVy/JP+3Cgpy89gKMU9NAYCYdr1pu9WrJWHATD3n0vQSLz8Hb6xVjp+nJlr8Vm
aRvH+ZxCYXAyJXcZsHxo8k2WjyQVXX7CWBgX0TcA+BBAWVu0FS2LVriFqlVaXNiM
L1yyrw4Ikd8RqP9I7mCFkP57FBhixoAgF8VKJh8SVtTjmRQnFrSJQjqYdWo2NRfT
0t1O0bfLwvMO+NgqcpwZnSL5AqWGLhpcB1/LhwSvNsvOf6E0F4RadaXSqQvMm8rI
zn0fNsA2X8usISQh05dLWqzrMsotjTzkoPrPfiHYdC03kCPQkfi3Q/yAbDV9n0CC
Bq+D120XTWZOFRgfzOMQfzCIPsKOZ8+Ntp6wdpC0FecNCECZ7KsHrjkdWD/2tQfv
3C6ojn2rNnq9WMn52x2vlMyKqvRK3AkkzLkkk37+Ssqf6DdGywC26Ell6MbnlRjT
d+dcRXVUWqy/D3n8HGcN+w==
`protect END_PROTECTED
