`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SYMT16tAriA90ct+j0nEnfuDBAGa1JRicR6UpuktAoQ6
Uu+Y+1w+lBd28CWqXehiZgUTvHbgsc4SiwtAaNm56Gp5n3Avo8KVMiwnQ4i6ShKd
5pd8dingw5Efke1SpW3DwTpBjHckzxH5jInpVmqrXs+/NgvkWwjlhBZTz6eHuQei
`protect END_PROTECTED
