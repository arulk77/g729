`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFeFlBvSdn6zLtyK6MObhDRB+i/aIvBFyDokfMuxFpmS
uTtwUA3yCmPxnjHDIeHG6qt2HOrp9HiuCYFTzSX7R6GWJl07noWQVgsY2+2gY1OW
iy1xuc1s+oBZg5PLH8pvat3NAkpzb8E+hUrIEWsUYDxCyuALP0HmnYwny4FTZtnc
I4EOOB7H7vX2gDcsMtvQgt++S0IZ/0dCbBEnSPHrtLAgP3NicimD38hGX0zbQf8r
Pk/X2N1dYhWfmrUSstAglynJNdxo9Y+1PXUZuiwMh2aSAL2rg7lYTajnTr2MuLD1
PcWvxYqDizgWs08xh+pARf+j/4WgvmQc4zkLNHocG9FpFjVwxgNyNjfWL75SGMvl
UpeGUhFV893EfbOy3h2gQQ==
`protect END_PROTECTED
