`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TyiSn4gQws4EtPgRlZljvZLCQpteuq313BEHkPsuGMyxGsU1eWrnwo8rXN9yP2L2
H6upQRZEYP8FYrrA2Dyy3EQPTryqjtnd4iU42v+qtIdmDRMn3sfbMJ1pCPDB3uY/
dWNZP0ffFkze4CC6wvz/N2HOOCyOscfyYTZObnxub9D95oiieh7M1h7YzdUmqLLA
`protect END_PROTECTED
