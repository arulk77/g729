`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMhV+KkO64ni14YEDTSPOAjtQAJBjdofsDEBvdS826ij
N/RjGzLxSpYBWSpHCaWEX0dvMzP7Syp0/iaRwv7Z0IDkiNMt0ScwNPgZbUOSGk5k
+hZOPq63kqFYQcQv07y8zJY0GpQ2A91InTlodW0xiS3LroF5rq1KDztlB/dW48nA
Cv9mxS2+iMlK18ElMZ5R8X+4BbVnbllqgpOnWWVi2v7pzaeBtAnZ7Drhg774cEfW
vrtviHOZnkY8Ojwx4nOv4Xb5Ux1bprmZUOC1O4WyjLycsAbUY0B5ijHTQ616Vjnq
cn2vj3pAUVBRc+dl4sf2EOpK6rXOsLmKE0rFUl5q2g3EIbNDWlCmNfNMmn3WXpuZ
t0raViOE7ujzilQpHKSORkYCrbbv46NqYM5uxBdk8alW7Z3YC/UE7nkdtNGH07mO
5nIt02xOPTsO8jdMffKAmuOPa9lWfMi4GVUfxX1+MSpHTHpLtnO7lABw6KhXuChD
XqNXHW44/YNA1RGxiZjB3C8jSGUSiwbk+eEAvqBP68MuSqed9yPvNDcmpFQdeyQS
m77LyksCHguLH34TZtzmym1nejcAhhQlNL4K8ZnwnWw=
`protect END_PROTECTED
