`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40LSAmyi2DJGPpipgNoDwsLv6P8KTmwKOIseJ7oeVPt2
29La3JVXX1x6eW6F9vnBIUUn9Fi/FSeep2ckmne2TV6PTMkadO8AHzMCJTTk8eXR
cKmgo/L7EjXDsUyu7m6ci1zgJXAFyJppngjPC7WBLRXx3CxFGGj3Ky8LxGIaXq+3
hRV9VUlESA57drvnFZXgYQvvlKL/ItpBD20tfC8TA9QopcKTIff/rrcy613qLa9r
ENkvs29s7ZCvGdw+ZPzDc2izva1YHNKgSzPbYc7/ftSKB/lvlGq7Of2vREav9eDH
LRxjhHDaEJLsrgnQXD8NLA==
`protect END_PROTECTED
