`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH06JIN8kljfblvMRcmOISX2dnze+/Z01xc264MnNwX1
uKPOcobuisn4cOeZmWT7oPbBnnigIzFJhWODwW+RX4IEy9z/RstV26zNyDb6/kYD
+AOSQTlUv3Jkcm7sh2yOc4cbaKhD1W9KUc8JXldU6j4b1k5kf0x8RmBtf/zrcYir
`protect END_PROTECTED
