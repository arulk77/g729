`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEL8ybc6uoTMlZgaIXxaqIlY+Z0p1BA9YswePj67LfvA
zGXT0JcnTF65cfA+cl6XxIGnzc4HT4z7gEhO1jnSadTst8RLDh3Ol8Pih2qJ/K5W
MAcsPj869BmgBYiviAC8l7MCr+A/rPZ/MlStEIVav0uVxIWv7IzzPO6xU/YP0V5V
pK67Wk1r0GJ02CQdTXqSG+0ULVJmlRRcVw607fiLc75gzQCbTEO9MHLZ5WeCApfc
TUn4QIMpW1O0EskjGr65gDWQum4fHkCE6fbN1zRtpvEbS0S0EqIl0neSUlBS1lry
aX/JuOe4acBvHBK73eFgtA==
`protect END_PROTECTED
