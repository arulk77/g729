`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
8Dmspv04ctxyr0qc8/3+XfaWKlTuo2dHhSvQPI0Pbxz54lstAEqkLeZVWweqrvEy
LQcgVSNV8yZcAI830ZAOOfGHI87lt/sxmE8HeEzB7BRrsPM+KyVGryTxlwdRfCNE
m2iTyLT4388h2qy4Qjh4i+uIYgdC6hPrv5J4wMT3K1Pc+HmyozfREhxvbJrcCMEg
fSUxoB3Qcpc1vpLr0gx+xDM6ueE6izVTMyd9gliM7REP7DBAotueNjUOd6eksbur
`protect END_PROTECTED
