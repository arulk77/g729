`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEVoRmiC07yVcYq1ITUr5DLSlkwEBzfm/daQJ5cxs6Rp
ImzKE7FYRL5HV5VsbkuLepj+uAtpDBdtGPjZGJx/oWJr1hm4hie2V5qwkUDLjyni
GLlYi9NXC842rTLdx9hAe46rmYcp3UfBUiOU5cJI5rR4fNwBrUdN88ufrT8I155y
Izil3xM4jZ45teAPWgxvdSYW3jIINbR4Z4yLtzW+ufec2+VyTXX9BsUgTT3AKauf
Lm533KDTq3GUF/h6Ol2ISO2IyC2Z6gOsuox0fQ3m2pfLzKxSKIeYCRuGEyHJLJLB
Bm29+OrM//YJ1rEG8Qs7pg==
`protect END_PROTECTED
