`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveASMHUlbli10K9ji+5sgfg2pwa2oaH38yRoFkFEVtyxK
B1+NvUqtCntTo22495zIdwmKKx+NzD46jJvnPrFtAGMexDpwI2TaDcwHaSSuMISn
dl/CeGKy/KTYhRi7p3CgDIHabtd8+nHDj3NxCVoYAHJ8fiaarXHupDH7QJNpi3Fl
gS30XWB4n2LClCbiHJtnmfwPgpAQuSR1p5CKVy2ycusLIhNgekJLNaHWbGb+gOLL
`protect END_PROTECTED
