`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePdiFagWhZ0HqRs2ESu2osjLSYG/SkYAqglLv6pKrjKG
w55WAGKzuLRb0jjYAvr+n5cXLqr+1uJey2ikfR47dCETydFtFTOHixugUV8DtxXx
TjilG7gGL/cBbWEI2pjVXCERau77Joy6J1ZQdK52fa3stFa4cIk7tDExu7ldubR5
FyBZ4IVLXZvAo8G9Mo7s9OQcaZx+tPLZCMSj6NW/WZTKdZ5g3APmbn7tt32ucx3t
p82zKgnAlbM8LvYzTFdI4tHeaSmLnJbx7bA1gV0wLReQ7lYc+CkZhJAfQbDTznVc
3TXfzm/ymf9Av4kIoiC+r4Dav+pZIBXq8Q5EohDTvlZnw6rvNm5Wq9RE+ouMvTb5
vZxXmOzVnMdtI/XciaNrHjf8WTScwZADMuvx5aOAU1lNaefNiHCUDJ+w0gy8NFmA
mK5tvpnssgbsRmI5dQdNmXM63v3NU9F+NhWxy6R7cZ72J1P2zAohQ5MaTYC3le2Y
FHDqwYt2bTFJ/s0i7JLca8jt0txnc89GRFtXHcLpy7sXpofo2hvxmnuDBKGwu/M2
sOvroS5fzq4FBWP/+2Y16onu0fnqLLmtFh3ZxzzEkA5qMF4avCbepYpALz2Kt5+N
PVvAqfXpB3PZHfKC6hZJdhOMgwvc1cCFBwJwGeGBNvQCcx3ZnHMPfr63+zd44sno
`protect END_PROTECTED
