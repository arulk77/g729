`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePxmvGSwc3W3nDK6lpklUrfLpde9sAK9uNHOElnFa2QB
3LU+R6vhYqAVEeeYTzL4o5oapQXwwWa6XPtzYn2ekbV+hQjZUS5Yxvbibpd3IAxq
NnQDxrmxINtwJu3x0TwY9H68aKyf9JTVjqWQIhBLGNSIU8/3vmvraYXujMVJCIAV
LnliRVsMsGBTxwyJiHQ+UpQ/I6SLlKNFzKO/8BXpAaCBUAuQPLq/q0TgG2onBty3
g/yMhxla4qqEA4Prrv3CR4nJ3KzLLlsUObELAAIM7PUHAkjfRM/A6BgPbwmaYKMU
qmygcv38Zabqra/hYzNJaiPmpyFXSj8Q4dpyW5tk9GuzaK5z9qVYcyaiJMRZnE7n
QWlk0hjLm0nAqPOEgrvEcqVpLeW2vy3SKU35wqe6Zqe1R5xpspO5jmBfRqRuq7Ik
Hg5IGIS4sLkA3UqBNL/uHFHmYXvsuRZcxODdNf9SMFwrLjLwUkkW67sqzhAY1wrL
9pzvXWE0PUe2YRCnSM1xZaiIlGRoulPlL7wHHLZNXkBHeFn0h+nn1I+mq5aW51AN
hQ7jRzFGoHt71br29SqjKDZcYvfggSSlJO4527dB1DWfE0OmJp/84PbvI2RTX0x6
MDcuGg+Mn+VowywBY6DbitPD9PP7enc9GXP3Ryl8qw5hAJxnn3nAXM93I0X6sOky
y9DOwiDLMDSjk+go6eOKWZ+96YcXBovF4pfPI3fYfWCvrZKatQdJoDBK+HInn8Yg
v/HD8KvcUGEKNC2BjJg+/RF0RNiACxzYTEpGgVbn9L9iM4t1l9aiSR9nNKMLbqcJ
iZakwh2yOhLqM+2JurcEd6Nizdhh4gYW3hYDSnGuHfw=
`protect END_PROTECTED
