`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDUezDuu5mSJHCuSoEB7sv9bEA3h+3qN5jnd4OC/u/2f
pEaDcOsCMeZ2BHpNHXH1zU+1vbvEWUiwL5cAOxJHLmrZ/+mx+tUvQT0FjqQA+9Fc
SWTxgCjx2WIkgHCCbRrSUGDN3hMc7omU3kl7OSImyoQLweArxtmvB5VzY9/bNb0K
HB+H3pNIGX3PEURV5kRBG6yfNZG7cylG3NJKaDrkc5h0Vvh36tDYHgFmRKiICBHO
pH6Y8OjW/FxE85BDKRsyBrhOqvkbGZZHg+v0WAFNX+dvWjPUc6fhftQyfHFhnSQl
imT+nZeeJjL5XsrEKChYVmbZxngq67N7ZxcYYOO0sQCmPasNJx/Wwq3+bFiGMEGo
gv21NLzCg4wuZtfdk35L69u79JJWdv3ofgtnYR3EN7MvgD+XrhucYgxKXw4pewyZ
/Fzmj1jCpuXV4ZILsiE4QndTtaONrID8kTzjo9SxOvOQpJLhmH/a1wgQaO4W9vIn
Wo2G+mhO5BjVSbsykRUgTGqIgLfRV+/aYaY2sIjsamfwkufxW28YPF9JMHnlMPiW
7egRLbnO7UequF9p+mprIuAUI6Hl6mSvjNEAT4Q5YI9NKDV0wE8qSm0zoADJO0bR
7R+pr6I9Iu/LbwDr1YIEEhhH9H9Vy1m4x8SovnCoAVT0izB+mYzqCbIHrk5PblRL
s5mx3OYqJ74EoGrtaTGGOg==
`protect END_PROTECTED
