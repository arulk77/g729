`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/MkW6a6VRx5PdpBbIIn0+QrfYN+d7pzGwIp/t4BonTP
Z3bfPuU1zdi8ZzpKparpFOijcBfFBbKGkGKMuqyELpPSQv5epq1GSRaPooamSm4v
6m99SnyEabiHn3Ydl0GJQbZsKS8VE/1FEOKnO8fe9OqicjyOnX+Qy5ngEYd9FSfD
Kk8urRenbGunOw09MkpnMePv1uCx09BMSy5ClII7Iv3kak98oagVr/x+vRGHiS/+
BheuAeWNrBW81VsMLxwwBWOrp9kY1zQi5P41IydReejecMzuATLSYnyUE+MXuVRl
IYVkEbbf6rrt5qsKnT87M7PAKqcuzxAuyIthAtoYFd5cII+T/YClx+urROPKuRWn
F12nTXmkFsI1D4qso/IrkQ==
`protect END_PROTECTED
