`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveId/5+SRDPkSmQeMi8WGzKH5RgugHVkXXp9OVexbpyM0
ioT66fdwmKy6bH+shzqQw/a7czttufXcf0Jaf0gTd/AkckNHQni+QEhEf9gBQYzx
9tHJVEt46+uAUVNgk72gakBETJ9qm1Ffvr92nZ4LaH9Xel9k+0Y5UGwlvH9t3Oos
/a1sxk7pCzUZ+hb2dUo7V993ziPSTYoyVGNTJhN2u168W+/Id7SSdTSvEukdvadf
bpSV+w3qSgvtqqTy6DE2dbT7AZxA8t0FqjFC7qk34bolECn3fCY3ol2BbFNSlY0n
`protect END_PROTECTED
