`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIxaAmdRNX+0hu3DrMxYbWbdMfApB9RWdGRbIUvMBZVq
TgFDXCbeMpSWbQIzvh/mkBujNm4WCmSeKKFu0UPwhkPOnuO4l+vDoGiyN1Hg5f7i
t8J1ZZKVH0yoyS74kux3IxUlFcz+zidnfpqwa3eMeUyfGk7NTrcZJabLw/um46ee
AC9zWQ7U7lu/toypWf7vLCzIrcbw874kHag705Jhkz3uPLh8pFDF2ZKRkQKJeWwQ
mT0JplUOjELv/wwS4rELnmTut1DybMq+GriOK5pgRswuDu/wKgi9FQtxODwiSuv1
Yee9i0DkWnJeB/dfrHEVIH8DTtRwhSOH+Mo+64Y5GWRwEpCg05QCD5OpTxK67N6/
+k8RLwxpwGyNbxjIJk/nZEX0qTOV7tqqxziS04D9oOnACGKJZmgfOTHtiApEArYB
3QvmOcKrY+YTszDyh8GLDopjEV7vhOON3SMy+AlXgV/CMdEgz/WkUslaE+vnxDmm
`protect END_PROTECTED
