`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOGnxlFh4ndJ2qhFcQniV7NstsAwRfmzGlm6+tGlAFI9
JqtoODfZ0HKtdlTUhPv2KvsSH5Zj3uHBLsznLRg1evXgo7P+NPF07iOQWqKZIu71
S+zzK8EXZ+C65Y+INMkvraHGI7u2hfq0ehFUo1p5qckRYANjeMeMw9+m1M6HI53t
UhTxyo+tNllVuX8wyW9fJyBf7ak1Fn+1vfGEdqA1xtxJmhn4zWYZQPE2EaEf7DvJ
iH5+ZXW+2jpVtYt4hY7ous+4ShecOV7DuDp/LA4/4C7YS+4sMXx2hkNOPBDajv07
euaaCichb+otpdaFt7NWClsyVLBpY60ADvE+TiJX+qDIDGSXSu1WS6k/zErD2epS
GCsgITw16X2gRCsnv1kC1A==
`protect END_PROTECTED
