`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBD7l37YyWiHllVCGMUhQy0mnqlQvmRlP9RkOMOUsmmo
i/HeKSJeMUPO+Rb2pBYcbZyUCB6vB1i8iF9z45o+9WXOPU3bcrKDgZdIGgspzyP+
UC0tJkfBJazHrSOsgZmEiUUVnBiOZhl85ubPcX2706+nT1BpVjZojDvQh55vFN01
wpAnJtwRlBQjxMWvyldY4hptL1xjADyNZcTKNULg79nX++n9yaoAtbUY+4U5oeGD
MVh+s1ujCG1XDBm+USYzmAjLNOGr7FSiXWIAitcajJZMJpAxObaapTd4JWJ54skR
8r8oRDqbD27gM3jNd69KuWaGtmB8gV0oOVmHLl6Led/jrVexC82sgBobHo1BkuLg
UGHYwqmqL/moA8RlgwoEKBriAymOj0h793AhjXcHO9mF31+i53YP5xpeGDpeLeYw
VjGGtvreLLGTHqaup7SJDGIrvV1kDjTGlc1vRzP8g2k2pJVp66zBqzIbiuDE9iLs
Z9uVNHVtovYjvldUg7MWsBS0OIneKkdGvgP7e7wDeXT+nLoW7CKqSVRPE/DPTh1z
`protect END_PROTECTED
