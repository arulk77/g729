`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOl8KAjIIVWRDv6FTfjj3sLgWgx4ySJGihbImD87sKb+
6T3mFhsnapEt1GbPxGF/OXsIPsHeUaUk4taUbmv/aJ2UOFMV9fLDnaFoRKw1WQfQ
/Bjl9EbYPJe+D2dI4rS1180ZKAGx1u/6XG2kO5o+v1htocvlfrdMWj9ZloV678UR
KPFU9QzfmpbizYO7HLYEg5H7sR3mWND4DBzovS75LzPC7X7qerA1yMMqGLeeqP7J
wHVY9HliTSJjlL0q3nysps7I1PTPv8LZotGGSUSpwkNEgI9LXLL7Mpb6LkAq+WDT
dzoJLxRsm4VV3aTktl8E/A82AY2I8SU20xPfR5bE/7Z8Ttsv4mbslPuaarbm423Q
JqWVi7kH69Er1C8t96HiihAnwS9r/RKa+jdjxCsD/AjZxb/2MIZGXuLCnH2Bd+A0
Kph+/y+S/ZWgWeY5FeoXdHKFsREtHq+aT2HzxyzlUDdAwsv/5jenJidHg3tj5nnh
USbShj+ypXrQczj6F2oyuF4gArmB/e0RK6+V4/j21W2MTHELJ4ZtZksJ3yKp6725
`protect END_PROTECTED
