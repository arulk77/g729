`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBZKifiII+taLG48SakvUcaOOnmxE96KI+SJIcb/Od4d
I7jeo3T7cl8Ai85T0p/E6fqWa5sQzw3OsBg6i7M4WO+m2+1U8P2v/CsWMaXHaWXT
aihwa8Bq7i/GXyd+0szQUuGEXfwmSM+FXD7A6XtqzOMwHjzSd1YhPlegvnyZpzZF
H/z9Fs5Y8yv6MHggbPwP9mDFnAylmV0jtdJgJcfH4N/XujHdcW1xz0q4W8/eLdsG
u3Eso0NBsVs/zuzlak58TgnYLVRhoJ2QqvcTbO5Z6cy0ol7mpG/q2QyFB0Gj4CYM
QBewzyb2aIxZmjFmVmGach24Np91hhqIJnOWTf4Hczk9jz0LtBRBJ7uRcqaDsSir
N9e/n0H6WAwa8qlcqAEGgCBOaYi00vvP20akX7H3op524gdWSM33lOpRa35L+u51
2UyXwl9pgqw61pYoAEmQT7Jq4ds4BZoEUUNgkDZ33JYB1BMKAhYDGPvCedyRh9Xf
EmRX7vLUvcW41N7P/hRYU0LeFnOw+7TqqZF0Zplu1tq2SUsZY82g3ACtsSgB5l8n
uja+XRsDdaWOBi3IaJJIs/mvGwveL7HrHWPhb3tqLsfZ1HuzMqK40XWxqiRfKUyZ
BxpYvDdojRbMif1wj58OlI2bLTme2Wj7YgANG95iRzWiYQEUsmXkUYAhz5gMnfJn
0bUggWYSzaIpXEwq3psQPbKC5Vu9t0I1fE10+LLnjukgGimChU2dfWpT9nDG0Ouf
6tuZbLJQQvPut6+EzGyF2qnSnkjOGGRaR6r3btaIDbk8xsAvux3zIk/7x7m74xce
RgqYWK1aTEBNCrfltde6XBDZ3gWtW3B04QuSRMRMocg=
`protect END_PROTECTED
