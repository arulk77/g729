`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKpKSkIheT4/8aRTZenAWPC1ow1B0Uw2reOW9DxImI+p
iJk1OayqotDrsl5tmNBvqswKYxeUg4Spoh+kvsIpTONXGVYTOIeL42h76xxAkad2
H+2uf4T4OpkmKDoepLOFVPq7NQFjvtGstgoqD0z/NJP+bwoLKgnhWrU/8W0+k2W6
x483wDzDO2ZUTfP7lXsYAA==
`protect END_PROTECTED
