`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHCGj73nFUm+ALePehtkHPFTjoRqz/ogDP9QuFeJ44Kx
cmUth3sBEo/Ih3LUtegXNWBFyAEVk9R2HeMFQMHunTJ+xPeurSHz2w+f7mGQHOxW
C2f5D/WcI8pOVkgG87OXbFtgui0EuY3VwUIOL4sMeaih6TmCOjWMR+nTCBiKSxPK
M+5yVZegD/vPqi6iDx5ktW9uxZ7FXBrmu0duWSTHwo3D/ZRgnfSKO7VpS0CaAIZC
vKo3mLfg3dlfioa81hcycXE9vJtZMl4I4VgikHD4vH4=
`protect END_PROTECTED
