`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJLcfwgYHNaipjSNfMxVYv/wFBv1cz+TbBx90qqoQjr+
FB/FMHtKn9OszXlZVhMkQa5B36wgCwI7ycEdbw9Cuk9+yijNe7FixbaPtbF/iKHP
CT3F0keWgZPnF2vWdETJFal4SF68NVlhbXnatGf4q/aUWhjdToVD1qOnSo3LKRT3
w1PFdDMzqIriPX5zyPd2Me/L9hYfP9NDa6oFCxDDvUWb1APOg0wY8aCJCblNhHm1
zLWAOup7JalZQIEx50eSe+Y9skFeF6859R8cgicqZZC0+7wZp8KVmOQvKx8W6DCW
Fbc3TEwtCeDp9gB0IsE1B51GGInO0mSiWiclLsRmdaN5IpfEXEglfGWmKo6Zti0S
Zncj4n+7vo/nSrpINmExGg==
`protect END_PROTECTED
