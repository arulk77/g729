`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDncKbvrxNEEuMZK8hIUNQI3tJaoXPc+kvDvsUqD/Gr+
HVyi54uR3RLPgJb/+lU3TryMkwEWXAGRU6QPkyp3TtAHI0DsxTvoyATzYytGniJq
74RoJolp4e2rgny5uS2gY35t5kdecP3Fy+TDWYaa8NhgmGbJl5TofL/w5ypCdbwK
jMDWTBznN0IPuipedA9c78PzfcKWsWP88Jnq4DgBK5hkVxbOcuOmmrLAD6NOxY7Z
jPIgF7vRZWV7T7gMtDDdSkrSAlovPREkrXOWI0St6PxHn+ZSryIKkf127KopSj8K
SMIxXGRHWk7u3eC9XuRysKKlJDGx1TfzEUA0OBkS0o3KyHr7gV//ayi0wRfbKXYF
kXdCHB8l3PKiwpBKXTK+CglFmDprcU8Sl2vriZihwzExDfUD2rzibsb63vSzOgGS
au/gkYB5bCibx9Poo4+dqQ==
`protect END_PROTECTED
