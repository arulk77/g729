`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEMWseUZ9w20z0rzNsSymcPE4S4Qr3zWKSFB9nAtu4Ks
Nv5cepnJDzLUb1VD+aH7FcRQLiNKfsArlM27C2A2IUuSj5Ukfc3QVUwfc9bzp6dV
3/RQussDdy6CwwrhqrnDoU3bX9a/lToD1/dXPysmZwiktLWAiSHQko3Cnag/aoAm
zFcFxhVEiH2GUnV/9yceKOPtKAZCsYhzHqEJhb4FAZYlJh8qy9W3F7CH7Stdu3uw
GuRf0sbFX0gjIWzs/0Epv2nxjq0P05+IdEwHJnbiwRmsoTqNB7lBtkOAqYRr4ps0
OIfx3IXJzbPRv/wPMJbv+Q==
`protect END_PROTECTED
