`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3ON6twM0bRyFDJLDX3Tyei64Fdi1W7hJnKQjvyu0yVSRRKfFUkoOrIh8D8mEDnBF
HH3WHduXM70bgHoHjSXi1G7XglCgP/jHDvEYIeNcVFvTVSSmseHTaoMKeVk8ef4l
CMdNfGHT+KvYZGJ74IIUurfcU2hrQB5HXD2Nt4CCukmc7avYW46sWQS4WRc2mhBU
ANOS5NoazS7SZh7cL1rtingyM6I7wX0XPrzg8etZ8DOzPuRsHgSYGhixUWjRy/Ow
W3Hn340EZTHxBC2VjKBq2VdCkJw0eAbBBBhIaB6C+J7vcYknos1tnP5qN3af4Y58
`protect END_PROTECTED
