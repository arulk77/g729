`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGYciOGIButPrVstMjj930qECMrFhbxePBlrQzfafyKp
8nTgM1dJG9Y5w3VARyP1bGf5eWhAif+oWJE39sJrH+PwPEiyEnrplHI0Ln0/7bm9
yIlxMuhfNGEKQTEnmRqAwl+O2sEPRW8S/numRfHdy4jFnQej/GgrrJUuFK8WiMWq
XS+YJHrVYDZS4ChW5yvoBg==
`protect END_PROTECTED
