`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLGkfGxMPGLpwFJ8bXbXe/IXdUgZ2Z7pxCwUC2s+2nE/
VZAuc2qvyxPiQfoj4yRM5eR8f9P//fmgZMkq0FLWW1ef7SDsSDpL1LgjDm9xaKUM
TFBI9G3RGhQhnicViBIvBtd3oC0PT53ZHzOQ/IN2FNWfbQDn+DOkKi3ZOEKag61Z
EbCwPzMtubkK/c0oOc+wi38Wvr2LBRAwcrngMFx8fdlbIl4pNLMpEPyJ+LEmuY9x
VvzW1Adthh/DZRfQ8zZU6lJq9J2cDcJzBRr7oZP9XfL5awTdIXAkTWFbXOjNKrqV
u397VY+E7vDqjULIfr3T3DcCS+83kos+IFONa3krCOML3z+8i/Y+0K1MfibvIrCa
t594BGm7M9jcSyUb8vyMQtt8mFABWEbD2/SfL9GOt2g12fyxZU6fJc2abBx2+aw3
GkFMS8VGhsFQCIph+hcLM68uBKbzFW40AGlzOY6HvYW/LgK6kguDaSOfo64unGlF
jmMGVp8SiLiBjbdSV6B/uLSqq/ldzoit4kQziX26gN/49VDKxDO0tiIi6Yuy/uBJ
`protect END_PROTECTED
