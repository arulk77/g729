`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mJp68YnwpMeUoWY2hmV7ZYZ7WC7ewWNKsbkL3YopGZFCEOuO+a5kHSExr4n/k4TV
UnCat2DJrQQW697jp4fL89GIAnjcWVNq9iWxen9AJPv2Cm3yp8VOl273jaKpNt0k
O/dmYYbFDTz7Anpr4df6GlqSD0HiSlmTgrTe+cXExOo7e5RT/m+NHTti72ZlapAg
1P+CmjXfOgcaUKkKGH8PwZzNz7UMNewiQy7816bsJOrck5//HdpL3oN7crOZcKfc
Ctq9i/qNV6bse0eoypxCzVk/xe31uNF+88dGcH/0pjJUfUiuLxLA+KTLt6G9zv2I
235wzu3BnRtboXrUASeV7Ca1wn3BOPgio9zGexFj1AShtO9tLTTNXR2zuxXMEVgy
yH2hyHZfbvrCDYmOwI3hCv80PoTU5PwVIwK+GqoiX88=
`protect END_PROTECTED
