`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIEX55yS2IQMjcn9hsjVTrpdCaCMKSyRTt47mc35TUtQ
CmXEwPjIzkFmigRoyoEBNAPfa1im8WGav1m2Dz4DF7HlSTqeR396+6LQPc5toRoj
zXQEB7GEmmfomAKP8ljgAjxW6oNGhVX5/wyY5nlNhfllD2JWH55oC7eEOLHl/H9d
Gu0lYh3ixJEXDfAXy3V7CSHwfHQcdfBWZfBGXcLQ95NHofiyR5OTNQ/dh9kBEnuf
U7sCnbRIB/JRdIxz/NMcvw==
`protect END_PROTECTED
