`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA/HdjH8j0rw5qs2/ZBKsa77mJbM9Jnjc4fy8UEGAs7z
vPwlnigcxD8/kqjTnEZv0M5glCGknYmiDymbWWy/2+SWwm+zlPT0fW+RmeTFmCxV
eaewCI5xeHnQkd0gd8koF5G9loxemcQeHVWrxhLoGPgTPpGPvA219znCoHP2QxQ3
HZKQjas0TYD2AbdBSBGi0sdRhFCcu3xBpBbFAOGB+Mu7KU55lMUW+MM/vhPN8ACH
`protect END_PROTECTED
