`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkTXVAle0xzfio0qI9JGVcHO+FWc+3oAXL9tAlde4H/Vr
zfR/xU+8WMTu2E669LhEd+OIe1AdXi2chwtaCyoN3D3GogksLNOmwFZBw9j3YCxR
FWnWpeosacNlldOzFz++wA8Jg8oE9x/RHAdUa+jEP+Z2bTWp8XNA1BtDG+j04ygQ
JFeYfmKIL/LkOgZpJbjnSbCujh9JJzv5d9Ok9flgYREJ4dNbGRuqaV9kCaubCVpY
gBRZB5zQYjSlY7XVZKhdHXFXBX3jCeEQcRRAHLqG4VTQin+8bi24DDEUtusGV/We
y1kDZ/xlWVGa9vtOqxHS2GdaqJl9ql5siIF4K0ivUaumbu2evE22GvEWVVm1wE8z
UXpojomKbaL2U9qTMEEvZkymtOVzqhH/hbzfUFqXCGM3hRVnXKYpiNnqiIl+dXLK
8VxwlbfrTsyr3FM1iQ3XChKbaL5RMik5Rdebu1nVanXU9kYxoBLl+c2aeVcbO4RK
ZQzY7oNA2MwiYCJ4NJclkZNFqn331pAjfgQKlyRqA7UDD0hi0i7gvZe4Y6VostW4
i0g3RORLG9rfKZVUA+WVepnpPRqdYiRt9S5yrJyYKR9FdN9WFeSD2A2hCb5aJBMx
Bbgd8b2zMSGQVkMuo1c98W9rNjhf+bvg9EtGYiNuObWxg3UAt1+LT4qQs2kAZsW6
hpt5orSlyBMPNOALLAygeV59FrIbXRH6HMaqsqLN9WuGBaffVE5lxwszJtxujuLD
os1SEJyEk3C2BWXIRZp/IzNbbOaSztf7HDA4+ewojaJrLWLGu0/IoMuXFSkgCpyU
LXznyjUA+SESeyK831IZKrSDYuIEFL+/R8K30j0ptLg=
`protect END_PROTECTED
