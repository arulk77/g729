`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu454tyHcHtT3A18N9iNB9opd+0qMhJM3PYcL6DL2/6bjL
QGJfBFw6q5yAEIwV1DVFTQB6lliHV7rwvp1ST18c8/tDv3L7j6TyfMWRlOM83Rfo
/Rju+P6QagK9mrC32NZADc3sovLHQZqqyggzpEPavvNRlSiHPTv+XlZxjhyjv2gN
XUS1leBimoR1ooVkJwWhPVCbF3YJRnyAJf9ci8vjMNzAX+uuS//MaQyqmW8FatZm
WTW7jBaYN6lKV6dD8K4qH+YokFhOHrD2Ir0GB5ozaTM=
`protect END_PROTECTED
