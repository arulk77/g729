`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDq5Oe+4SS3zRZQ31kkaDYaYmDsTHhF+hXhrBbk/1AIJPR
OJzkCC/mdm+LQBpJuUuEPTvSLI3ejsciHrP0y2608o60qO4J9r+Zr/PFZ9vc5oFG
upwVMxxyKrXu/06AohUtAgR0Ev5k/uYPCP6Xmcs/yEt6cE5E5YTNGqwuJAFUBCJO
zFrS/jSN2kHONy5LOJQB/hp+jPYQ+bwTh1EH4Xr3lVGWXPVu+Pw0ccPmJyCyA6wy
2Eqn9c3Au/aY9akG0kalydawvlGtH7puMsCczirGU5lZSrKvKDkKCGznyTl3O/kU
`protect END_PROTECTED
