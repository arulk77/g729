`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN4PKEUxKYrWQITINGyW1+jsv9Sz1nMxW9ASrjYAGWT9
OjSIOLFWtKOYl/9H70NYjbaZE5d1nVu7SBi8/e3mLxK2YIyzjgKOQRjnmoJjJ33g
K7ZLQFlYpbZePGTOFO+Kp+pDR6cQ9NUGOWRslFFk+e6w+Uu/Pl+We/lBBPl4TDj+
WdHhP9s8xAqdSntjdo14jtCtYxV/EfyqrATduKTWTcVdf/MoxU5zS51DgLbGmdXz
ROCo95neOYIItRxslgJrmCoTCe/ot6v1xOKNTa6MvTE98OtA/wZXMRaSK4ok1eP6
i2Z5XF8L5Irn2W2TqOMt6Dscr/yM1UERvOs97guauwdoyP6PBaV4Jv+MfMKpwwVt
DACiMIF4417FOyrBvPyCMgxdcUnKPEw7mTUtoUZ3Xu8kYC3GvjidM4uXG2ds6LZj
7t5FDHi/v6ehmQbpLogjV8T+hsZLmYmc9Al+nlevT+qJMYVXEMV7Im4KT8OUNizJ
cK6l7yC21wR1TwtkOMw3HPBnWtJ9G29Z39nvYkvxOvVED/g1IR0UzOENMJJqLajw
XV43rsn6KSBDKJALNxm71+uZ8C+1R9wD5mfd8QAN6hE=
`protect END_PROTECTED
