`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45bmS8dKERVjFjQqJo7nk/O0RnNgVZ6R0W6k2YUHGkV2
aDV9QH0r06tjew0dYeXNzFcnDmv/TiqgumTK/ofJGkKgbHhxZuvjkKU10ixFR5/Y
ytPlKD/Q6CtVyoImpJcf4ZlwdLNB2YLMQM2NZRR22FfSQlm4pyQmaItkBWdhNOw3
lItvB9tUJL68hv2Uh2DledkLTPEb9Tu9X7Jp4HggKvJ8GgR2Z8P2zHqG2k9rxcvc
3dF2KJkUsf9Dj+AM2q+xUGfsXc9IAQoJAxBn5ohjsQyAFAqdle642t3pHA4mJ/gO
YLfBFuVw9qD1DO9oaX8vEQ==
`protect END_PROTECTED
