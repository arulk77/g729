`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
05i6+TZXhEozUMR8mpvI7d0uchJzWri9OdXXgBzLjZVLn5UgEyQ4s6bEhB6o+jmr
IeOxvFY2RGU4fojWkgBrbcGASz6gpv4JcBUAq8lBN0y99OorqgvO7XWAEccq2tJQ
wyFfO3phRVFZJnRgk+x9RFxgcg0aXDwQeK6MKZLjsUvJgMdn1RPVFemJOxSerVoB
zbTFKhzT60FGWNo7oOvRWYHVVqLWqy4seU13OWhCmBF1cJvxdCYDvNRB/uGYjlrE
mrmrLJK8DapFqmIu77KRlHD9DK/84e2sxEw1WLCrFc3waousw7sJYuc+gH/+eSCI
grwSEFcujjMumIMBLnzmOcl9Orcv9eyDyuPnssI/GiiwASH8L35fMDro4GWWY0zP
1+Ditb5dkofNfzHyMOZBKrXa3Wq5qChYtiHiAJLoPIgxSS11bxOtNlkwxWQ/PiYt
vLtelmiGXp2XLhAdSjSIWKvlZkc24hf24n09cVbutPnsl2xL9As+H8hUlYiIP1C/
wvZwxYTh9LHjGt1OZOiaUOt+iUB3bOVBtIIpzTZTcj6inlF4w19qmgJyCaSxtKJi
3Nuq+woLSaxLU+SvO/Ts3G648nByq5HUCYrC+G+bqKImCvJZuum+DSTm4RepFEJi
ILNEAEXoyUmWnxpvXH34k1IUl7lFp1/uZvVkZ4i3JV5t/K6lLGDYFDuzNRdU2kxw
Ko/kCcKxzQklF9s2JbIZMRAeUhyVKLcn+5qooFQli1kUbDzZqYpC3vK8JVWsVlKH
KP+j4XuI+cSK1yN/OmaPJlARwfUQ86cyIioZK8McejnFV5ZHnIAQ7lRZJjziMHUl
e0GEJfnnyxINCYCJkrxpF1/A7ikZW6Wh0Y9iCaENXdIrsrgaG4EYu3B5J1ONAHam
DVm8kpQ1TxU7UFtEeyyo/xiw9yDZT2v6gEqh8IrISjk0VdDMrQoV1dn+WvZknlwp
cgq5ui1sD2AoMfi+yg/ejJ7+/MMY8q+JGJvVDepOdmvmEIJazboAgCMHfu2JbJmZ
Sd4fIFL0h3sznJ/xgYgrH2qsO6x/EaIsYqzxJd0/UK9kuVFKyJEvncmxM+9Eo1XP
vEXxIKkBdA+VsMhluwLnJUjuMDMay6WoF8Jxh1oykUjl2gIGfuFNq0IiZl27SS45
GzVQAq6tmSYI3mcF79sheOuVu1DlwBJ1prgx1YBubOqvfY2pGHMUIjxKeB7QqaZr
RXqr1Q5M+gtjIDV7pD3OXp10W4W8In9Ucccd9vPzrTU=
`protect END_PROTECTED
