`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f7/abUqhjDM5o1RFuBftj5Thf+Hgs/803otKlWIAzS9ZvoHC6B9rJpfy1Bq8wjTf
laMGp31/AXBhQ6QqQY4n/4frUxr39jr39GnXyDZsLoUvBwI4XrsEiJzqlYQL3GMg
2eykxRbJg03AVYnttXUT6aY/WnGAB2OgDc9EM0w0ybEDBHGr6V77v1rDyBwAvIoi
zphJwXM/Rjgam4ZVMwlG13+IjWSJ3iResMobNlLMi6TZMTzaPutkovqs5F1X1qqQ
Ki4slgMtwwRjmHNxYIUVN5HHD2cfhguPHEFHR7H9PJrt/zDMQ7E6NknXrL5PAIpT
y9cnZLu+xiKyTa+G4CvWMYSyrZTGIeght1as2CAOb8ufeqMqQynd3P6wY/4vso1Z
Xu+zj1vvoLm7mS0F816zLbstfu8B4arvY9xOY+oN9a/PAipqwOsurESPjGYCiCO2
WIOxrhjWL2jjg/Td2K0y9Q==
`protect END_PROTECTED
