`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iJUbFmMvQpqW9d3mgdsysiypnTT7yocqkz58uDD6LPa+8fHTSCSjuCSJLIM0ve0M
bUhi0H6II34y294GhoakAQ012qCoGTYX71s/X/4ia+yapxBwzac1cREaB8Zt5a4R
q2S+Yp8Q/9fzJBY+UmXMIL9+l4oO8B3zvkc2QOyByu2BQj+ls16TpyAY3c0S6h0c
FvCX9p+Spoi2N4HxEOAVbw+f5aHzevR6+KV/E1Wb587VjPFIQkJyEjKv5julL2s9
jtDPEJhzi64fwZexchtet6yBRpJ4tRDZKThkHh07xbhOZD3EB0Wdhf02YBQQKi7y
9oX7n/caBS14gjR+LLx7AtrSob36E6lu+/uPX/za5cOC6vzuyF3CGXG1qo+GgBTS
U2MBNKS0gm+pHk6TUAWru0ybYVgKLBGvcESuuywBTLSZz+Q6WR1oYOKn3VT0ll0d
csmeyVOnG3bXhjXyH1wuOrZvHPG36jtQpLC64oQk0J2QzutB5FC0EUqYY7Yh8cWu
XWxAi0s2XcWFggVN8p2MFylqgge6H2/In0+s9CPT+nRBiQ7eXUqa8c39h4mTsS9S
uJ7CrVHAotGfqaiactOahRMvDnlJsSVg24Keu4IgNQhbOQt2vs6zxpRyou9G+pmS
p7Y3cRV5GTWJfuK9E8nUIZV7fIjrnPP7pgHfOR9zpax7mZeCqsSMeqKkSjZvSMBk
tULSgCeXI3fIfqnNThD6PTz2LTXd55hsu/7OrPu9GyoXrb5+fRUPUyqMQ9nnsgbZ
a6e2XC41v5h2wgmj7AxBGfDyzYDSlsoHOZAbFaucDUP2gjvGUI7Sqf3M5wqgev6c
th951RI4jxur3jx5LeuSx+hp9vur/FVJJ82f9MOm7GA=
`protect END_PROTECTED
