`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GXu3xX6zxQSGrM6FyhZR0qcmo2t17kApO7OkYgu4PGS+qtWKyH0XxpAnbYdPAWje
25vJeuIuqMbjU+jlfwr07qtDvrkE2lPizORopv9synr2W+apOab41FuKmBL1C/8P
qaTFy31zaIAy9emnGbIxsGHgKGxq6w24fXlXz5Voo/JFiJrKFvgEh4I4ftMgj/dp
b99u/uKAwxs7IDvbMu2Iu1oXE8G0gejDVVnXbc+tyOf1N9Q24dCcR5w79YlmojhT
`protect END_PROTECTED
