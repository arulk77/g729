`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAe2XsNhmC18QPOYlXOWji4O7GssCIVExPC3qzhBVCwT5
8KeVcEQL+g4KXLTC4sStajqweB/RNQtf0dUhApbEmEExDXsTcO25pUOWn+pg7Cna
UC1CozYuX4TL5aJvVG36hw2oMTWL+K/KiNNE1xDYPdP7dGxLpZtJrrXJQ75RCUir
ZaaZuMrV9JC83ufui1DNNuyP3DMgzeBtyX9LJXzJkZvSvVQ5Fj4WhtLQkRuw2X+k
nfpA/zwmAnfGTFXj89nbQAvqYI4rIjwZT2tzxIjyKXAlqMveMuOTnWTN8kPIpfLu
Vv9nFGmjuSo+IZYe+DJZF6M2vXpJkFXnc8j11LAfvhDNFfq5vwMme2qlsMD1fbQG
VQKrIgRktfabdRKsdhiMVIWqfvIIshq51jp+xB6vpUJ0xYEmfN9VMIIggWvhV/YF
PK+Z5mJ+W/mWDtY+y2e3nFShBME1s8zD3rFQx7qbs2zNHf4LAXeh0nBke1MVETWu
rzD8NA7NYCzjROs8AEeKsrvZhi9PKygbalWTCbAS1DiACPhxQ6W3qkPnZM7Jwvn2
31+pZRwdO4QlpdUBvyDs8iZw52iePKWLVYgrDHrpc5CP69b6F/NBd4Gki9eWEifa
OMJxcFEYGmeGQ6ubW5QRVJFs8Vm6JDilLbikaYQpZEdaZl7wnr38b/hPMxnj2Wra
5gN+MGYIl+VRcE0/dH/eFjaydXo2rflbnJn4TfDBq6hs9P2vqOXpKqV8mgnUWNyw
+RutB1pmi1zZLGk7gPc+/xlzSocD8GQxJONJ/H5PcwTG8Ok3UDJhe4AJL4NWhWRg
8Yai7B1y3VQb0AoIpxiWcKQkCBq3ysBs7uGdvokdTkms0n4RkUr9uJlbBXiJHDSe
EZuBQ2Pdb/jurUanCnENMOzNP/Zz/q0t7BgPnOQ19Dw7J3ecwaSd7+RDAL9vWFwT
0xN6LdoLKynaHRkC8JRR6+hASF3kBsc6yrHbUNFHET5oGhedN/sCMEjE3ZXxLcF5
Et3TWQfPIhAONqf423y+qG1zHlMiSSun6uaHn77nSN5cZOuRwaR9YqWm9UQMByrC
wnmBFL0JIie5klNI6AkvtY5lKhLDV7OsiYKk7HJ2cVfxz8eyHEbDQXNPiVRVcm4n
jTVjRLqM2WZMpvmOCYcnBpjzNRaAcr91vATxPtZgYEYM0YYBcNKvZhxEic7oqlZ3
7dc/Ak0SIOYRKiI+sGj1vVFXbzUo4tqOlgLiLdZl/BDqptmptuknYOefWKlyDvVy
ecGnc6Tm+mOp457eJIq2PsoQCT6rJqOiLnm5qKgx1lq+hP/bkpZG5czFZmi+4fus
6+N1E5mdMGMPJh42GK84GoPjooHpplwumEsryzqXf6YWjd3tB3j5miXzsXFa9zG+
K0USAxXJ0GvFK+y7Z0T1Hg==
`protect END_PROTECTED
