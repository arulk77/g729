`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3tIUFzyPnI95ic+DkvUUGqDMR4yLQjOlKydlt6CI7Cl
1UE3VFm1OtlG9UVRT7G2jGtVISD0k9FOcr1Jm/M73UYoS7nZ1MtMaJJaXs3ZscTO
OzCrFXIN/ZDffOm14ReaT8cFsOqUyhwAh6GBSONVbQawKiPX2bOmoXEoi177DteA
bgI+HaFjktOT+Me7nq02fd+YdId2Y1PDH7tcXdzViO/Ph4Xvm54/wPZo1vHO5ItL
Poez8xEYowXtzWro1Sf997zR655OygUfkUJFmsYu0sX9hSHOtGEWKQebrS4Tr1il
2f1rjnDPLFLh9SwxIrmyMvjJSBm4Mi7sE5gKrh8jntwWh9P76s+nVVr/sa4Cpagn
zrZ05cKzYLOo7ij/snq4Dub+qoi7thRTqNBeKEkw6EeKF1IAmlF584lCZT+2qPnr
YHutQH/OSxdrzQyR16HU3pUdi++lxHE0Qp3/9T2zSJNt9xQAKyE644XNxKCv3tZc
YAZNX4zM31YDE7jUOxh84qQrY981q+Cd4pdtxcZwV0GKSYhflEfHTAtRL+Ubt1nx
JoNwq9j3D1dXfV67xIf+LPu8ZDwcDfL4nMdMgPifbtbYkvBx5y9bxEhEzb2uXeVs
mXghX9xkWvgBDAIf3bPRppVENHJToe5gfdhS4VPIR4w3zcp2lOwBVgvBOUiwkt3E
scJSSHEwy7KNDy9D1O6GzQAZqKuy+3tVd9q5jTuB6fdHgURg2RINGSddroN2d506
0Cwj20k2MrSmkCMG/YLGcoIiR4jla6cIVFYeXeu+xq+SQhX7DcGpWRRSZuDQbNjn
Tvi844RWKCj7XbijdavWBtjJqxIjgvfuYg4uTNn0yD/dxKZxjuo3hjX1NT6sCQ68
NNCpTmzfUqiLOLabYsh0s9RzTH2kkfdIzPY0pO+E1Sa+wAgKhPhuomunBo5eEh1g
LHWdDVHCZIQQr/a+4F64Q832OkCSbs7lehetO6o7ja2pGLPgOYT9mv1Yiryz4z5L
ep94SUg/IIf9pTVkUqWsbrcqKX2CxaiqnBtxmp6u8fh3nYWPQWlePe6jnBYvkcPN
1gCNk0I9noFQIjcnkwlVriUUBuP7hWje/DJASl6f4OB8SCHLu6Mmw7lXXYlXDk2o
9r9MCYbhI+TtsJcASzJeIaQmZWkM8weeYvmkllLAdJayWKVu3SasuOsYzj9zrbSB
07uVqtAhjhXm/1DwidrM30zS5iaO4fYRJ9Y3jnj6XX8EDTPx3XHLlAng+S8Xiukp
qkkVgLYEzN3tekG+7gGXvwHK6WB7Qg6FtZ2T2kgSKid7CmN9EkLYPTl/1Avmgbus
ygJCsc0ys4nPBPXDg4VWC5zH56zvoVgsy6jPc21zSjnrGdfKjUUp/xaGTu3kEF4/
WD7ZYWN0iggGHQ7jxrlRvcScY8TYyhOIgn73UqhZt2WfvnGl/wguDUqwmN5W9KYl
Z5wMOIJ/qBphgdHe/Mkt3O4FiKQ+PlbaM9NzeM5v6osVLeGoEosWhdwsfL0MiAO5
ryx/Fta+AQ9+CZ1pdR5cEssOPcW2cGtDfvPM2RouhnAZdgb9qX3/j6qVryUTNrzL
6VwEPF9l+UanpJ5cSMtjJqKxV8HYERyZ80jgfhtOJ0vva/QI9LQXbEA+ZJaYhrHf
MGA24iR0E69rbOj5XbzQ9QkJz3EhumESRkmqdOXX3Lhg3BaXF9vekn9DDQR1+4K6
OhblOlIQ1dw7d3HpA/fpgsDurEV9/TLMzpr0G31BJ6QCAtqYqzDC/PshR8BLjxpm
8qjcI9cwieLewf/n5zEay9GNmd7OF2OqSkdzFx2IavORfN7bbD3F6t/avX+WqW2K
E2ODczG833yoNIfc4CkmNINxfuQVuy3y0ts1hKOexYLJKNnRvV7d4/D8yJlkWR5W
sVVAj/nryqRNW/zjebAqMX6MXlTIhdlVTn8LFhXMUlO4SjxXLage8Xk6IswZtlOp
05aWFXohawXkWBJ5pivHdxJNJLMj/ONM0Ql0CEgH+5Ka6ooFenKcn5FdtJhjwoT9
u+8YftCDzNkf+Tk9tlX04nPJdhBF4QFD1bADADrSamruidgN2QW/JwjnaA/A4qWX
XhpwKvyEJIXbA19atDkl/lniGpDbmyu/N7OQxml5HhYy3anQFuhCSMDGuQMJsUcA
tp1DxO/VI7MaBXEhhxWy1q7pm8zFXnI9Y4qVq1ysLo6k2/+Afybg4v36i6G/5bRy
U8KROUsXjAir2VKE3ga/hZvd+/DoA7KyWn2/HlSWwTHjp5c4b1I3bHwOIdxNz8DS
F0+iEmbs/EXwh+ETUy5jAqgwnKlHC14UpMC8GnNSuw5u8jDKValVk7Ah7ON6q1mu
V51KV8tzteQWgkynueSuI7bPy/3aUo31WmUGPFyprwbLrZ5LnNd3zuuB8YGPT9Ht
t6+i2GtLo+kmYK3lCMdzuP045ZAUGx9ALmKMemLPc5KnLzm5UXIu09S0Rm0xpzrJ
QWbprA15mlub0nwv1n8aVzQPMm6ufltzwebzsao0FzCqGkj/z7T0m02S2C4bCu8v
EYU/1R14S4Sn1e5u51M/razVDGhpXM2l+3Sm/6vAb6KvoEXGucvw8q1s8bAWrDF4
WijYJHZ6BcAuF0ijBrrsl4/GCX48/GHsTKCVbe9Vuh8eeu2zQXAeJN63jiIFMom2
i2JEWalpQ2N3SwJ1YWuKtSa3LtWsvg2QMYikCJ4SDmAwV859tsoUHpjP9M+tnvTv
VQ5SWgvpjQUenLKx+mBSirsDo1CXCVeFmQCYFCji+SBnWxSd8hlUiscR6d86c1zD
Xcju1++AMUKpGVQto7YMWcmJsG5MJggkfb3RxxhuAAliFc41hnGbMGzNb2DjhpqL
znUc2wugrdMhm/viLut159nccRdoHTjpvVqTE4mf1IvhkceMHip5SpZoHd1Ty88g
6hH566HBaxtJAndKV5WYUmRu3IeXM8tTR3UQFfGMLLwDf64wkrznhuM0hH9PNK6x
bSpNSzaISQ7xyAlCnLNE2fPv6wtvnRo8jP9dnH0sdKBFIglIjUUHC5QaeAAxmar7
ziVbFzhVmlZHlPHRCQqxIiYtjygh6HKB/EclaftskTj5pzMfsJ9/xoY2HOpu7ZC9
pSTA96P7cOFAj8gp/ypSdzRIJwgheqHHNITVXqqWOby6GC6aEMYZ6apuFEDaqsjd
kyGpX4NutpENJP9itzRg9VS7sLr28i4h7geZzspxbh+3ah2AnXqXrWtmDcuol7/p
8Ya2XfElVRCnMa4M5Aj+GwKOPjE1Tr8wVCcTVnJVtVstoKqM2wlyAwRKOd1T/LI/
52Ah8h5bw+mafrC7ThSa8MV/xUpzt0CNSEwWSSgLZUw5Vy7DrHkarAm1m9pg/ozj
GuUeEfgiYoyyy+NSsTbvq+jBvYG9Rzr/OkQOr5VCcQNE70jLPdHhvS9HVN+Kjm/Y
vXdokQ5NYOMJSKdVqkvHXp8Oslxry3d8lAeNhIq8BxYM/UtMmNGfvVPO/wQuaUfu
n5nX7W7d6BG8VaF00UvSfWbP46Npyc3YF5fINDp/M3p9vjKC9cZfMEx1+9dt0Q7F
lExA6hoALlBl1QLhNtVG/HMtGUWxbDcrdHG+FAZU832RpCZmdb64F/M1GCIpAl3W
I+YX/fRwM6Te+E85Ig2gzkM9XwWljU/Q958GR4Nuise7FDIm0M8GKZ9AS2dUJU8m
awac1StBqNTV93EaU8wTn4OSL7emB6wq8aToTy8j0zqcEYcL5oZK61x/h2i8AOVO
2CD7QAdlTV0AK5gkvQygwMA81/Fe6/MrUpcFiQULQMa1PpApx82pUBA3ey3/j9/Q
TjRz4Sz6KnAANCQYLm7Bkwxvyu8egqenL22yiWsaqFPlVk3GZYc5wUhIAwrIaJlT
DFtc2rx3MjESR5LdJX1hyOMqZSoKZ+Nf5y/BXLVVJRq5f4tJAc9K9x8vekbmcPH3
+jais9nc4/byZrOrD+53NN90fwYJ09OOlvhdIRqDWpRx8VPj/tMzpixBsNJMYRi2
xMqaccW50vz39UTFybxVzYTGdV7+0XE4G97Sj2dBd1YemKJru4eG+5u9ghauu1Xz
b/1m3USTSETAQN+KJLvMgCjXQg25KXkATXOwdTdHtQxIxmvKmU8U95NOSwoN8pBD
q+SXXjgRXneGSW7m+8pHwJ5P3IKnvD1SSd3U0HfyeJjlUyVVckAZAkPGjypwD1Zi
sDu1lqSmC3+TgBDuxkmyFtENxrZIM7G8SJmYxOiNkhxStFqgDTX6LE2MSwWM5MZa
RMtqtNgPy5k65ZuFS6LrCrugq8OF4nEy2wlr20apI8rqhuXEeP/+3hE9o7lkcXjG
HYlM4Tx4aN66V7mdWzEUCERThaIG96SbPMW2YOmXEDHzws1OEBLnkYjf3OdaXr0T
HIKwRhg/Uiet66u9KHq2BNcl34lHyYhdCHgMbvIK8l2yCjJy5poPj5AKgH9GIu5+
4PaWYWj1YY31MrsePw9HxTD+nS0vhauxPxLHcD3/TDq9UTdfBWWq2oY0Fe9cRTl4
3rCkkXZRbNNkNHGWVdOzTBQokA+kbAZ0daKsqzaY2QRPJ4j2T3nhQoQ0JgAVdxw0
PEeYRinPOi4xanOtOvLqykbIR5tBxaH97BzZ0LuxCEqInlFtRbWmtp8aYjY64gVY
QhIn9cvMFgfDS3iqlWVvGsmLFrs+B2DOBqjQ8a7zJvsQACdZIgkdxke4+zYgmGZC
/tVPi2av2UZ3/hWeZQ47rzgA+kEgSrrkc9zI6x2kblItJ3wOnkNePemJ0caAFVk6
HE1m1AbRCLN9CEG230kvN0fjSqEvDr8ZgjiwIQbJmhQfWB/Wt4LPFunaqVMkqBD3
U26ZncRdtXvwg0zpPRx2hNARrWqiX0r01cVfwUGA7l6DOsnQ8GFNnfY5GFL47cQI
wEC+ZME3qdBow7leJdM6YE316g42uPKMZ7kA1n9dMUUwzv/37xOxvgwAtJ3/6pqL
3y+emep/tVzzCS4jDeN7MaHhgExz/NG3foRlKToTBOIZRhWm7MSx7eOcoQFBdNPK
ofiaBQNN7x3qwefQoebPPkg5hW7nfb+5qzMywcvp83Rp5fKMJuPBABzxeRItohWS
fWoBOPXCdPEmL1XGlRbeokRDw20rLGgwdvhZmUewEPQAeIs+227sjZ+5q3mYGAc+
4tDcDf6YgqwL32jSny4zMXClGGLhqs8p8Bw9/jBJ7JB+GkIK+sR1/jlguPXyNVT0
SmX/Ec0ClLPJsiNHxKO2J2G81hL/0vYqIfK/ckYpQ7NxxALJO69GJsCf1QU+QL9A
opHYo03E4c+MEwpIP/M9qBtGKo2S8R0aRCJD82TMwi9duodBjW6eUu9X2NYi4JEg
E1dAaBhqocHH0gcKIi137K0FRSen200wo25/RUPtILgm9ddyxUsIi4OfvTvEc943
H6S2BtnCLpuZr9N/yrCS6cbv4ZflqNX+H4dbb1+uJc5j/JzdwGV/oCiDWQ9osQOJ
8M8U5laXp6iIP2gK8ZWBZkMqc6ntQ/yuRmu4b7+eveTBsu6rU9KaQQ13pSRLC1Y9
/OgGDOuN/4i0+m2zOhUbew6c3zQxXtAohVK9NkzXS2hyiVpSRaySL//HYFaHricF
9+odi6T++kHE2RmnT/TgQGYnqYMQPvZx4j3Q9XhYy/CY50CJyS1oPxvdFOMG+tkg
BPPridrO90yi6L3qfbQUJlH+eqphIduHBiu7KPB2LjtjxnAPW1LGHItfzzabqwDh
CtniJxHaXoA0N9XXrVKRSEAvUx3wTtesuaAQCe9RwXJmRUYm7qaErXxp+LOjUkKq
Rw3V8SGKJIPxv6KU6VjQFNKNcOCJjuUnFPzatB4cfIlZlOHkHiajp+F9umi8l7VF
sqYOjXsxcAmBb5c9n6W2F4D9L978evcaMvX7S/UUiTlZ3lDCTp/P40jdtptAkvVZ
8bJ2d0EW9X5ULtWr6G9l3nS93FWOn0OhpyqT1/fM5ZH15iTdegb+4PS5IXnGD+js
CwMSui2taIURA/hG49YrMy95wCJvlJp03fgZZL53Cayrr2K7WHIKjmoVZjcTrDDx
rLnwlUYscjwhVQzeQtolC1eqo1H8yGHMoLyEHszqGu4Jt/K5reHjXReNUpu3qVrh
QBhbTm2J3L8JM21TdfAacHWbaD68V386HP7OQEoKnQlplSi+L7uTvEISpl0zF2Hd
hK2XS2I01F1CM5nVCWP8+2WanQnx+W3047fiIVdqMOmuws9qVeG0qbHHbqLIY6DY
Pzn5MuSZh/7PAkLW0WR1kTa8AThGf90yT4aVJSTmMnZAApWT0C9yiwdLTuI5+JA9
Q975mMIiyJnAbTI+TibD50NIgzqUpkqqLOyv18qvTpLuAO6faiSAL7XaJsmPa1u9
g3UXVK28Au91eOiAzXX0Gqk3iKTwRLd9ziAWyfcugMIMFy8JkGJPdIkE+50o2wT2
kvAD66PayE1zu3SLrGKKDfBFQZXTn099HPHQMxiMa96uU/mGUTDExXmjpOQra6T+
pVsMcmbUoUyt99U/Hya1o0G9SLzXoZIib+BsosKePbleClRXAE7W1oyz1zxk0nBP
fyEMPoLkYQV9DSYDnQvaNyNp6WdnTuqLuxxABPkZ8dme8BojGUlfuK42khDsOddr
dqZmqh6Mhw2tpgdYLE1RYCf8BR8DqZjElreK9BAS/3mhwfRl7jR5tTzuleKYWvkd
1TtIY9a/AaggxZjIn29lIy7kf2mJXr9MCa6o7fT9o/4TqMlq5dg9070CKQAQkAjV
nw0aiZnUcxMDO9jLUNq64n0usFplm94bbal/rpET88jPCJQblZch6fe3FzbJdFQo
4hFVMyJDdjhkHAxfjb/YZOoY2YAB8J4MUrwakX/G6HWqW86lqYUKYswh6i7Qvp2j
kkpSv/QWamZUqan4dSSBHQ2diBxzJ3sg2BjpuULVv7RZyrqQO0F221w06gZgtR9A
WjTgNHsbvZhbgPsIXq+TqIVxWq5C8x7V/ioh6FrJban3gLZXADM3p73Xn26A/SRE
fcXCmxQpi286Mb6p9CUCzSgj20mpThOzdcMtnD/vze/fnNdtdIg1QAmfAYUFNsZu
h4Nlqi5ukrIfgPKGk6mnxza6vkJ8PxdRIrrsQAE6o+YCTzToRJUlOVlOf9swOr/V
KLPkr5N1hsc70F+BPaX+QxP3MuJ+P16RTbxbxThtLuMRTYf/ogjiWOePHM85odup
VfxLtCHwz4cQNXCAF3klP7l2Dp9v4hy4uasJNQmF80LL3natgZdlrJkXr5UtBQ/3
OmuVDn7gkmnNa1h/bSv90ugt6g+aY+6x9awOX1bANEjqlnJXXp8D3JwtDAufQTMM
Taw+/Lanz4XU9yOtSNopo3Vm4tgy63U7MznScjvKJIX2VB4aqnJZu5jmSjHLTLLT
01rSaFdN79sASq224sXLXTmqDUpndpvls6qRIqry32kFbPn3a9TEeJgDunk/Jlek
ZQitkPiubX+3EATPqta8CP1dGa1R99jJP6+6nYWMIB19eZuZVJSOcRZ/BjfBgmvj
obXGP93oBOHRSlgBE4xYEwrcanYvT4wbcbInOKLR72reX25Y4XaofZdkilf+9W0X
`protect END_PROTECTED
