`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bwaCb3ftkNVZrKHMxzXB4hokIQFckJve61lIDDTPN8KZlM7b1BkpcRaQydogE3SO
BEMG92HvbgfTzN2Qajww2kbCMTWoub0uyFb5L0xj3nI1N9xzAXjRlmfH5pXLAMKQ
29OCROhXwyZrWrn0odV+g5TdcQ6JZ3Fd3R9NYPiqWQY=
`protect END_PROTECTED
