`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePOh2L29zSNi909EPIxZ5/cnkHGSlT94xlho17qBpgNd
ZfTU2/l4zgcxlMOW73dVlyG9yHpzUEZCav+YvLvWdD4Zmn73CQcrvhrshgndsxt7
1QT5PQxfhduy8Fq/lo+MPZpaC9cGllozmhjl1WFeZPHmhF6lEchDdUe5G8aXsnCL
J/QdKvZ9qIylqF5X8MK7ed6HQKoVQLACEgePIoTX34LTggppdXYDy3mzK/ofmsnX
8lA1wmzBUwByTtnFEu2SWb2Lrj5GlgLCTFV22dcTkAPbPyDWk712mnCtuoPVZHw2
B+Z1ntC/exVaLD2StjlHvekef89vxb27kASD4xGJTodD901vxN1yDLrO55SsDkE/
1zMWa1drsQO7SdJ+JKh214xtdBN/PsPQThGOeaO+FR03gMVj5tP+Sr8bFkLZL6UZ
JJJTk8SAEQh6Nq4ATb3A7kqIJ4MtjXIRhMUvwtlvymUhrbyKRT2R6D0omvUKneaX
b4RSKwGptMDfrNCmKrTD1cPqtlwueM4HkyDO21Xj7B44giBVJN8U8Kq8Ir0UAFVu
7ItFF5x/XmeY+4pYpDdt2VVLvc9oAAlSkhRdoPZezaJySFMj+r/FP9ZmuUv5nmhn
X6JCAguhqou0b80e3IvzaeP+tBIVe9j5srhS+VeExuC9/QKD9ucL/7xr0ALLQ/gA
kU1qtf0czi/S7wPHfyOIctjt+WHRYudrJTWqJ265Fs7STz85PffUIX0dBSX7hdfa
oQEmuGTYg0FamC+/RK4HVif3ykmaHPhHiNg4Zal9LKuY4Vsmn5UGdYqAOD4FWqLs
nKSinGcJhuw6Ntk5pC3CVPmgFeo4N/5qNSCoS7Hx09fXNC3s6L6/a0GaU1H/DXQs
qc3Ivs3M0kXH6eYyw0ai0Bx7V1YnJdbWymnKOtKkTbK8jm5XTnUJ5uyWwn0O17wE
`protect END_PROTECTED
