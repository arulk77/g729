`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fz18j8l+Kpmakf712ziwHA6F8g0auXjQQiffbfNdyCank7WPmgw37Oq6OCZS/v55
mxpE5An2hFGtN9IKi468EWZ4XbubqK27w7fYYWqiSI8CReV+KbUN+9orHB1Qvbfj
bslAP4/DuO0omo8+kUy7k2LZWNqgWcFBV/vFupXV4OcQHPdScwg+Lh/PP4mlUUM0
9u5czWHsqsv/dlWCcdshubDp6ilWk6uuoWUpzjDxAtsM3XDmmu1HjUBrtm+kxQ25
e/CyGUA8R6ovA/zDJI757/WPFTaZw5KK6etXtV3AgupxnS6qfu1vQQh7CDnjcFW6
PPtsXTmFv1yFRwIMp+qWhwkJWn1TNRHblo03y+VZiWCDYoT3dV3SuhlshYnRadML
9+4nd+w7wPFLJ8ebxuhFgFQtKW9WATLa6eyoOijVKbFZLfQnBrKtT8jjbjzwl/6m
iG/YiiwMDg96g2osFsk0Q5SoLM0I+/U3S1aWl3rNnvb3RM/nAWT6dHY3IzR2DfGS
1DuFagf4fXSVM57X07R6oBNjqufMKLHOEYbJa1ZNiq3Cgwi5JrrKtvoOnhv6V4H9
bObny4/tBjzBvE1NuMbtQNs23KsVKYhl45woFGNEwDk=
`protect END_PROTECTED
