`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OPSR7lzhaRF1DxpetLu2+fihB1PNYxGAzQsOm8mqrc3MXI30N3xar8JceCkcT5w3
rbTGN1WIAczzeOuAf526vZGk69hiR+k4dNx68fdMr0YNKGUq/pa9ZY2zPfQD0LEe
Z2r7OVJfnPe4rG157aubpXe8OStV4rEGTfstpsYa1+PJOPBsa+V/OXkDRu4tCzF9
v36rQ0Tz3r5JFuKL3EpsevS64InEflH6ANwGqqqxY7bfbfrQCdwrtGtXAKN6lLaK
TfyHs32zyqBxbzZhLFcSfY7TOtvQjUnYG1gq6ZdlfGJvD+BxDw6WTSydFs7SzQb7
RdPZlpoaOThDicd2gvtqbF5dvfbfbsmMsIVIo3rVMiU=
`protect END_PROTECTED
