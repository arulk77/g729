`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ4V/EKpdiPyYQpnaHnxmxFw9NasqGrQrkQbkbn86Um/
jpthE6fOkl1vuUsnW7Qro9xqvrmrkCjwQy5oEHNAsymeyyUiDXMVtTvxbloP7Ot0
kATcgiNOLFhtfPEZbWET8MxNS0OKQcHysfN7HFVn5KjwuxxeaCBu4CehfS7r/ry6
vxXC8tAAircWMmwA+BuAn7fLGecLfvRTU/VKZsmSpHAs5Fp/2241EijAbiS8gIxk
UAPSY+Y9Ewp9faLTNOUMdJjFkver0+aIHohcHbRab4XNk7+1F9runNorJj0VAt/t
80YUbsbRPl0D5aTx2oPZb8YBbhl5cxMKO1Jt4RXIcWtMdfpQ2bcmvwPGjQB95LY6
Jzv1UoEN7b262OoYWvFTo+fpC9g8PbFBioz/inuqnI0SqS+k4KiqgENM1ZpTh/af
2/3Ev0bysc2eZNNQuBzA/Qx1f/Q8ClCwW2JwYJQ1GR1mjVFZGgBmAzDc34y9x/04
F3ZBwo63ApURza2gZDyyTSNb42ToYYH1rDe/tIg4p5phYGlSrmErCurozZZOoNkW
Qu7/Vlg4VXRkEBpgWll6G5a9FlCXCW2GyDq8h38kMc5DQxdEJGC6gh84P9JEJymh
ruLbdn62AugaH1/AwPXRopStsJCBTzU11cmKHjPEmljXMvk+o1NxcF24j2uNOQri
K5ZbzT4aJQTwWN5XHDXtwnhf/cPXbMg17KEyjlyYJe+TngyfcSSm7gI7PMlHY3ld
5RjTXJh63WHzOhYn7zMcplVC7AP9TEVDjTPA77s78Fi8s9B9FteYPnDGfncYbVKj
CyM4roM5l9FRXH2fhe69vcHSUDcR/XZhIylLpn4OzdQ=
`protect END_PROTECTED
