`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD7gKRRgS0Dhz/E6crGp4XrPmyWzkrBhFFoh48ZY7gXl
fDt5J5p9Vdmx7RmEaH7SDsasMwzKjYb6p06qRJ/6lWxp9aRazoOlgJrrwtENt7c1
5xSi1riX2jjN9Hk9gVJ+XDu12g8nPzrOK/woQT+UscgGGU9xVIRwsIgneEV18DYG
Rn6WAjLBb/S1aYwuGo+PaUltmQKKaEml+XZ4xlpEel2ezWUysblBp0BqliUVNC+0
KLcHdXpuaXkPsiBYQSEMXX2xVdGTAXc8FQyzrQc5y0t4o+yJlQzU0lrv0N2gcGN5
ufpPBq2/6gC43zWxgyWA/3NSHed/b1UyKlZnYN0/DddqvvEnPdREqIS4KWlFOzKR
KLJI+5T7sAV1UnJmle4PHrnrLzIHPDr8btfyBbrWi9C78uMVV9kkrGJn5+zlQnGV
uJXevZH+X57IiBUT/NYyd8gq3tEHkHjyktL8pnRdTzehNlri5PH62X7GAgHUzyB+
p5O/8GUDyT1dreWJcFr44x4YPSUdL0a9s8wJOa23dXfCNpPdbNPNHsx9TAUy36vr
b52e//o++AO+WBP+PoLPl/rVhJrtJwmOefv5Y14YCAYJUsZDM+6QoidqI5R7HZTJ
c8drWkV1ypXYGbMDlEbhonqaVqh0RvU76cYBVRMphNFpbvARuuHQ0xi+voexhLus
RT+2bEDeFWVx115+1nqNqQx7n/szdrUjxb9EIFNA5iDvITWjmUvJmaFMbgp9si3i
`protect END_PROTECTED
