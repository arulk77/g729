`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44FVbLTtJapJ2Mprm20Q5ZzzFFTysbB8W4RE+yqjJVkQ
aEk2iNvKLEQMWXFFVu5f/RKEoJOej4bHFZx46i3Lbb3IfGEmTqU9PGrArVhyuv0Y
gsiuOJPDpji3ODwuyVUBk5OYgqciOJU5xSR61boCPQV4yvPGH8Dr5HNaQ+w/zFEY
QU9MoflnHHcGBRb0PO8zyeWfeZ9VApvG0eUoN3ldpyJJP3aaoU2mvxwvt31467bH
psQruXRzuZRLosIOIbLfge4+Jg2JkRZTDZcRCVZTAWeuIs1Oi+yM9p0QFD7xB9p8
lriXiJuBj1PogFETNcnXtw==
`protect END_PROTECTED
