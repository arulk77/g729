`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
E5DTV6SflGbz8bNfjpbS3jBb6wgFHrSJjK8LMqiRBZ4dBGQLUNgqRhpVca7+Ktoo
oqDgBOEls8+Idp82PrxW2bedhsh5dOpRbO/+GyJTxP26nmsTUPAyD81XdThtZVGB
0QryiaMByIGSfbU/zUsZU8JlwY8gR1s3V8WDPRui0blW12w6M6Q9IY22Io18Tw8E
OgN/FdIILwhcdEWAky0l42tHRHCUqFx/3niV7o2JRtEQS+FBQBcoXYmLlw8B+b0w
KWQZSUY749fs+HMDAuFlo3lFSAu7DUIWHi84Vm/sMGw=
`protect END_PROTECTED
