`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNztAy/w5nWBBwGKcgHVMuLsGQh2T7PkheIWJKV8IGKzy
cd9byU/4SKE5km5blNOLJZ7FE7I/SvVJ7/SHkh35mlsNHauxGHTrgTGAuPz6rUNP
QpBa9Ywsf0c7S/vECK/stBmtxd44NlJNOfY6tj/rnJzOR7Bfs1qpmR615EwB0WVz
XH/CH9BSxMUuFYAydpwmRzQbT2qLYQuz38scDM5p9ycocYEJcBxc/N3S3FnqPwHY
kKswPlc7/yWrcPEmTj6ccauQQ4+WDhOrrhF3MY0KpIK1tgZGuiFFxxUkA3W5DiJq
2A7nyy8hPEQGXkIa0yJjJUr0q1702ZLPGXWG/GbZzVhGllhHRLYSkSDSQS9Ikbtr
1iaIeV906lJ3NZU0a521yEB1pNMCwzQq/gTbq0RXNxOH0U/L99sTfCqK8tp/0ek7
gM4TdND4/SGkuJHlc+aZozOUlCgOwMMXZS9sv+NHd/0kcumZFMAFawUiFbYhs5b/
0T1pWGeTqLmiN/fSOqz0YZmlsxUVJ8T8V99/3VMASBziJGBiWkCPmqXA7y3cAFJw
QQPYHYWLwtqsmCev9j275nWrOpianZGlIqppft1l+jHp8EjE2H9PP+dme8BiawBH
NTSPc400Wfr3+duvVclASd/F8jiOX22xf1NdnxDe6IMJQ64ymqqyTfpJABAni4++
sFnmA5yAKuw2cD2Jk5U6H0oajFY90ELsnMHwunbmKxMiOZ5JSTJqzC9yj1Ju+ODP
2D7+5h3qRp/s0XsQ7PvKlxPCYtNGCb64++drypxmWSc9NZYEUjG4Foj4ywydZKk4
gEiJHn++Z4ngL9xL2g4sEBvowhMDccXwI9nzfaLcI1b5RzpLJOA0T/B2PNKTgL0K
V4zrZcTGUTVVkhzd+1qYgncouOKU5mdEkkB+w9msR/tQ0vmYiah7Za8qeatRZKmM
4rT4s9sER/aHLHsqD8ZAz2RnvqwEfpu0fl2TVK3YejlgbD3qA6JawQ/vIZ66YLMe
Tvl3Haj3eF+gNOSjpdUpKnyRECX1ohNVaCvOHtcvvRHb8VL8jxMVnRcLs1G1Tn+m
O0cw9Bp0RVT10FOoqr01QkeKL7650hPU4Y66WBJjPycLFcWza9MK2t2i4cpE+8pD
YwCt1EibkfGeOfRp9yqqleBz3xILlxhp1Q0uMZDyyra6aeG6a2TbbelreOpXUSFl
ZyJ9lfmbHJUkm9RVCegpYO3B9yPg1H+tNHjaGDjeZsODBCr/QFrUWrwwaoF1jus1
f3BDl3P2/7nLA4r9hdVzBxnBjIBCy203/PCHx49vA6OAndqXtavYvUNws/kRyeH2
PkltLSM5rwq17KHHSTHryoEQbJcPPGfvEDUwjgXLozijnKyp/MvzIli2ePPyCAlT
8wG7C6cZ2hx0H4ACMn1C1HceXrkcEa147LoECghnm8cM7W8ZB+OneGXcwt0Ar4hd
fKMQ/HedX/K3FNJ+6vSy5MGi3VLIho0HwoZ75Cq1Nf4=
`protect END_PROTECTED
