`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDtuRICSiv/+W/la5aQ7kFHqQStdQYGrAAIku2bFK1SK
iNeW4RoRTmFDd5bDhvdv1UurV2LUkZbgrTfC3m5eD7d1W1USNLh3wo6z67zEcYDd
A75gXwYQWjBxaPPgRoRGOx7Uw3y6pHqVlyd6uU6dLadkkr4vmH0ZvjW/wSfZTvyS
EzVZwKWeBneMf9L8q/LhjHeSyt6CTSPrzFRs8wG4/5dJEzGQJCYBZ0x305glvOmF
PwZA+YG5lft9cHWXgIEKUJbWsIpwSwVrLb4VXkN7AFISDKORDMPf6bOylGc8uxlK
JcUa3TTuwpxHEWjc7E9vXvE7ABEb4rjyN+6dDFwADZC+IY27IkZFLxaeMgIWQVMK
/rkGseZvJuLWX+TB/ZGLog==
`protect END_PROTECTED
