`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5Kp8FsTBKCCa9b2kWYdk60LC/0/73PIuJ09wlw+soUF
Rje7r9kOF7GVppgPduviumcv0YtsgSzVAOSfYkbocJcD58AfzVI6fMrkaAfa4x9x
kKXjf+c97X3uxZ+BFCZqNA+BYAey+0qRl7er9DTorkI0klkcJOclSkUyB6Ay7sk9
LVS8+m0kfa4n9v+UDCpu42PSpIk1JIYviSNVYhXQAyf7PeB6NSXfYfJd7GTelmQu
Re5tAVGOeHCRSRYhPZZ+wTPdtnyRzK8+0k7WeguaIEtH0GiwWh3DJ1CChAByNOM3
Nbnnx1lazLLE2J9p9AYlabaHse7w9iNuF3U7gfjqlcjbn/ky/6D0OeWIb1toqkkD
8I6NK4KK4oaLZzWnUdPWY5JxDwaFaxdzUSq34FmAW8piv2/2XHDWsrMUoCmsFM/d
COydlK9uimB/G3GbIuONGblOA/++7xDm0BmGiItvxp0bBe2P/xsLacMqnnZb10tK
zdDrBBVix0rO8+FBXeqWu/iXukzzQdk1uIgbXETeJuzNreDnqEtEQo9kZpY1+lMW
R3JVwpCDQv9GX6iDad9Rw+vf8qFXKphXHkdnoqXhLd40ZKve35o2tSqjsUSB0Wao
fecVEbTCl/riIx8yk3ZtpPyzVR1Mq5jL0iFMPqDLpUKTtn4pFNLP6fvuOdC8EsUe
p5NfWaEG/Puw97jbfKeH2G2ftgS8MSPeo0NQ/7MQsI/QxumD1hafCayurtLnfunU
pTPWs5xTnP1GSoeFmFBj8JMFSTrYswy8fVOAWJ6ZjHZsrV1iuOjuVkkDBH13JOK5
IQATlSWcel9BewHSlliVZq8BsvbDuyovwNHtrRhgGJBN+72qeoDQbDhVIJL5XPzV
wuKSfKDjI9aMZc5MKgfFtdlv/YTfXUPq2cNquAuBlJAY6YZruqCrRAka1C5X3Q/D
PTEetu1ek4s1AQ6wKRKL53CKxQM+ysa+mJhqxGoYOE0iJ+9GUdNvpErDXVzQ7+hK
ySdHhzvfIJGPm/xWmrVc5M1EBGSqPyMVc3Xak5yNdStJZlsWtsqxq8fuy9SnR/fk
6IFCFOQhvsqffW9xoqqjYWzgHO7OvdjSRx8mwajL41opYCQ89vNMneEUigQcSBKV
NLNAtVGw/h8XhbhOcTkakxOWxRk1OuBOYmCFpueBPh04ChSr+gIYN4iUojLlpuHB
oE2GORue4/IiLXUQg+y/n/AEhh+HwHp5iYvCk53u24mgqSqh5+CQHHvV45JdtfYC
a97lVuVcI1ENdr2vDFWxvh+4U+E+d7SyBATszj3gJzvJ4Kt3NaAK5tocSZQy79Oy
L0XaKqg45hJiZDTiv/s2T9/Eo20IwuUwPKbMqApPuP95/XvPxzz8IGHypkQVGxk9
NoOoj7Ou46b6zm5EsPyrpP6EAOFO3MM1vLJlNh004Y92bMxeariqUKJgll9mgITx
KZFvMiB18DEDhXkvGZHOV7f/6xhCh2iAlpaSz7yU52oSYgIXZetNScOEyVeYUQHe
QYXxP+v8PZRbHFraaB1EDI3xj2/AQ5osKYjVtO14PU3rro1qH1Agh3z71HjAddol
NM3IN4DSK5JqjIH4NrAbKqa/kE84omjO3cUfGWFjfpQKFNvZ72i8wWwsl719QE3C
F+7GKW2ZARIjfYExDESzMpKZ9fr3kBg7cJIFnTtDHoAisex1hReyMNZnIjvOVlSX
2JsPZNtmZwR13rGyG2fs7bsnTq93++0hfcpfY34lDQcCfX9hU3o6pq9TLvP0C4sZ
t3zun+TMyoNubEBEXWV5E7X0I77Z94pT4uv2Mb0h/4M/GfR8jvVsO8Z/Xr4VsQfE
a3baMgth1ci2ogHRvckeOzoL9kA5vmtJwTSLpRh9DI2QOmIj0+a6Aqzn/I7zhJoD
vUlPnuzpCQpUubXJ6jvbA/b2Jtcclh411xFLb6gPGb762oJ2zQG5Up1kaai3IhAy
wgwz6M+SqHVJs3J1/WqK7XTGDVEQI0BkN4OAHG7p3F6IPob9B1NoSJPjO6jfLOo6
yxE4lYPi3UIzrO+4zbhG+znXmfeB01cFxHCUoSocOZpEpfoRzUhXSGxFt+ZArmEC
tAC0HZBcOsWPiNK29j1EQP1Tg3Gm/Smbtnm0TGrL9kaGcSiIZZLe242qa3YzCoKL
Khghw3uNYo+CcsLTI4lcjYs7nxYdcz06uWQaUNbXt5/4qUg32HLmQaTa0T61QT7Q
Lm60hsMnn3HQpydf1IeTuYtJvCYmhI+rCrZlQ0z9cwpQr0n7Hpv6Ji2oRzURy6w6
R63oNMbbrUCYUtP0/qW1tfBTB/aF3Yvo06WlnAR535whqCnrSxJJ9xmLJSYhGtc6
GxogGbN0XfGVd/fS7/X08esXBSv8ztdSeWK0Hu7gfAmrGIH+sZn/stUnpGKIEFnz
ujWgagsWb/rdc4KCtwd4LDz6+6tBvP6kvFOn7TKTKLOesL2WoxhtpZVn4uYT+nPK
O5OEWoPe+nmzpMYB9tG7tAdQ0H0okPf+a1aELtUPUZSdRgae5fpXO1xPk0U4zIwL
yo9fGwdRSAOQ6qfQ76So5sL9URn6/7qDg3NZQoidr2Cf3RUDOUWedYRDPjG23MeK
HyWCoQkTwWx518UUjsBGY4QbPwuJDYFnC/vVqqg5oE4KwAiyDMgsEbpLmOvveaT3
uzBqZmnqjNaR/GU2xrZBOp9HjfBPz1dCQttXt8XNYyxxsNetXsYbhLg4elx7y+KX
7USDYxhLApqufmSGkgBQ8iEl13HBkcZjqjXPUh6ReHBzc9gU9BRoauTnGibMv7GP
rdNOl0G0kjJLzqoXpBOCU7Vcb7vzJlpsyMiT1eFaEQO+wMRQFTrXCvUg1O7VBLoK
AGB1aheNPDU0uJ8/rlc535X9iUjb5WosVrA+a2jpECUzh1+e0IE+QXnCysi5HxkQ
A5EhsQJ2ll96arcOYLkoKSjGzOgT+Wqy9Pi4fjBpvvhcigVCsZGcDc0XYq6x2sa2
jo/RvR9833S/rLAc3jGT3UPVSWxC4DHISgu85SekR1590o2oqDM4U/4bBGwHuTQ2
UqAijWx6NHkymwGJxgEcZlEhoOuib3oVD9M7BYjOBxkvD7RaK8TiiTbGsgp1iL3L
tmoFP4QLRlZMs+GZv41uVshiglyqiFABM7M3lDUQhNPbKog6nrVmM4hl8Zbsr1yZ
bbmkhrDcSEqX7n2ZCnzzVkmfA0C/Dq4DH8V2xiOZVUwj0YPVjaZlPlHaa/CBhpQp
ozmKqY869Ztpqsuk0F3kjDFW1jfuH62OTeA9dWnEQCF0ud2gJRbcA92LXi5rZcz1
F5ygBw9Po1QG3W0hSUIFSA+MyexfBGZjOM0xWTlYGl+HTvMlI+DlqVuDsi59BpXs
4X8Ncv2E4jNh47elL9/ajojFQNIIh7Dn9Xv8Jn6yfgSLnDzN77Nrsp1FzO9PcnGV
PmEIdV8Hv/hgzGQLkSyNxrtJOCjsK9IL3K8QVOysCrS1Q4oBLjCtHPy9SvyGTgpV
4Xh06AK6y1UYcWF29swqSsz3f3+I+fgxHs1xsBiZMztFZshpSWcWijv2Mfz9Thnr
4AFV3YyftjiA11P6GuXIO5440G+zafP/TokHVJrd5J7qCECtNs9vxUma5dTS0D8A
xfS2HIxgmb2MnaBJ1oe537zfMr3iotFOdaJdtW0XAKuUv5U/VjPAAc5QYJDjz7gS
`protect END_PROTECTED
