`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJvwyqlNFcn4GoN01Py2Yv91dGjaqHA87jRPTy6ADg6E
aaBdiVcAGrKtU3rmTWMHcckF4/FPlETCnbHJciu6M5rzXPxavC2+eL4ba5/fN/va
iaNNxBr19pX+kass2xTDspy9+fg3AW1V96KgBq8LOOnVFe6ipzFxYxqQ5dQeMC50
4AzUH4Fm9m/ou41dsU4KhVxDZa+RGKWEs5JJthRKgofT7x9pWwJyfPsilItg6FEt
ytjj0s7BmydREv2+wueNsa0IOR7viULfNhr+IoVBf33fp+cjwuja4YP2wekr9npE
SjMRTA6YUBgRNWDaL2Z8OP1riIpeBWRiwknCDzNAFT7VF2cQucWbuQFGs8FzHSV9
eeOBrb6vMnA5Z4hIHnai7I5m5JXVrdcNverjKPzhW3b9/bJKOm6/nBbl4D/nreCI
8uMJm6L+6zjlWi8kvpD/ZeQHZIusI2sSfTKglOmPIgnxr80lyChthMzhMxJp0d2i
rwtKFzJbpQHjGAM7GExAggg0u+HtqhlHhAax2ipL9zgoCbLLMLKBbwq7zW7h4CEc
`protect END_PROTECTED
