`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C5B3FfQuBp9TkodYneeDB7YK5/TiOiA0Fg/gUYqg5z8Q
fN783++ekdpbyIbpz0fKndcccaYm+YmEx/lbK4PxPEiLyeJaehgEml3fhvoT9c5n
STGEz39Ckoer1jy8x/yWp4DrZ8RlxFO58yGpM6ZjqmgBOaie5anBFSorggRJwFwX
TpYlGo0bYEqPXW0Zt94XdlmqYW+StlIVRXoUO+IxHNt/gKuoJJCI3JbZd8R+JUrq
BNGxWAwcSmeVsmM83F+/MYJVHM0PjjL2S6lA+m98x7kxDpz9ZGOP0mSaRkya1U76
n19xpFSXhimq8q6rkvC6HvXix1R1AQM0CTZoPWxbjSDgPBSA+jIuNEJ1KLCi0/tZ
1DAk0KdP+Pi9U9ziNJtdOv/sbSQsg8MrUvzzEqjODRr0Rk0fzQQF3j0Ap1eTRBd+
Pj+TqsoIK0VDqnu3+RLBeDiDJpZhDfOlavwXs34NgJmw3hgLpBWZ1C+Oi9bw6Q0G
ua/T+m2wonEnrZ7qZNmRzIFDCzbGIgRbyaePgPRd2zHCxMrLpbXnpupyD04IpXzv
AVK05kYlcwB7EfOTxxQgr0bzdi9vIZrPxmzJSLOhHJEt5ND4jv8A15ztVyXHNMRr
rSllvhHDVQngiuNJHHRlJRKcRyvoilKe+zCdAn8a/pCdNtD/0+0xZtZKxN/gYFwg
wyoo2qssxLuz95WKc5O25n4m6ZvEnlzgnu231j7H7qxrIQ26A5vkbI9t0cyHVzGE
OtjGp90oIWUxr266LxcYmpxV2ocd5BNt81OtlWuq5OOFu7pDzjv7caJPgrpOUDCl
dj9k5rtu+DaMm+/Trej69lsFK027GS0fYKx+2wyMT84BQoFjzB2dfRqoDYXTeNJt
2cFnXOpXTMFV3HsDKQpTB0s5s8hUN10YVLIG13hGECg6ESaRTqhv6cb14rx5eHX+
EL1rGhwe6c6FclBB4lgWw7gO2AOdDgwzriiPHv70tje8RuLEBiayOt+okrT+D5C0
oMfBPYXmgdNQKyaCyNQC6qphRNClOvvpSuMmlh7rrXAK9WR4MK9kRIQl8VnO063c
DIOX/7i88zSac/TaVk07ptZrouLQoDT2qKtpQyefTVD48XksftsUOQo9P38QiNH1
QdeRpEKkrMyczrmhMIpeJASBsUaQpc9AckMmpHnKhkac+poFbwR4wvCVk409uyF7
iuTq6B7ye8yxnbzox29vhgYLLv85zVR7JXKr8WNJ7KgJFf9ebLAJgUzcESB4vdnp
ZphSn6NNYSsszjEpJsFfc+sl8DOiCMlJREVsfHvsGNfcc4ZaBlIMKbkyJ4+3Xwzk
qN74SXVpdUv0sC84OGYOonpUPDT0/V9u91xYl0qHW+169NfjG5aqnloVWbukJwYY
8q36BKaHhfWyIbqV4ZdUtJBEOxnaGHQKio8Txgx8CvcVIJAQPQZT26AG2kp8/lav
vuPKZ1h6UlMT1FBDnq4IYwIQ3w+JhW8guRtdoBn1cIoVvvPPx3Clbgep3lRXjuCt
VG3C1O+9Z8AK6FuGVWpwCiMVcNMf/9cBRNty7RL4ZfpjB5RSKXl2U7lOWHNuc46F
2pl0WBJGcB46HpdlRUojDRrI4BzJ6JKU9rkpYIBjyQSq3u4LUtpU+KUBNMuBlylY
9m//U8orGxdwPaBRQ351Em1BKrLd3WvSbdlx1gEl2XN4IZB0bp8zWpA6ehMgUPUz
OxB2s6bU8UV1AcRsBOQPjrqN2xsGEkwP+IyamjIA/amiYqc/FbIG/IgfRyZ0D68L
mjlOPm8Xfbq8RXIF1WWtIjbNI4iKvCEpxXsnBMkfvv/JDfbeey2ksa78PW+Lldx+
FDPStvyhwbyMLIbY/2j4IbrXRYIJbDF1pOq7CPePBf07iVJFwGuZRjbW3Q7jhxyc
OnMOZcKvrqfigLa9BmuC9q4U8ifbm1tev1cHRHPgeoCycon0p/PC55VppfIR6xiU
cF/VXrtLb1UPaedkCY/RTyJKLw7Jve8Y59dpZiHhkCDArgyvaRD8Ezb2AvdafswE
mGXAoj1wWM1goInTo4uTbSZbdR4snnWtRGzrq6pF26r4Eo/a0cv6/HfYPJVsLh+W
wU8NIoMmWZgDEGPPP/Zd6fWH3oqgh7QbfLFluEO/bA2HRiQXmn+0itC+RyPulYfm
55H/P8w6fbSVKDbkoMaXqNZR2oFmNK2+cewzJtNFUXY2aRCVlXbboKN2rgvYiq70
GG8RU6UJsSwUedMjExJJ/3E74Xd+E6Chh8N70K/UsL2fnkoqbCZWhEHnmUC0FygQ
sVRldiOgkpFHmb4V7UetajpvFj7bDMMcKNfgZLGMX6J/Rz4mlNDI9q/RIq9fNn4H
2+vCTmMDQbK1m90YC6keMwv7fn2ggz2mn1kYhxy66671CmhhqOn9HZwcCTtlrj+G
04jCStncj1gC9mqee1geQdSQqZ98W0f9tjkuTFW254Dyk1llyjAiqKHcyEUeCwAJ
cfJvSV48vmokfLiphS27TyWIHRfIlpH7slMWBMnroDADC6VkIWql8Ap7WTP5f+hX
mB5j6ZVH9hfkye0TR95PmWIRST9HYxXTPnnDMKYy01A416qRBh6WJ5rnuej9L+fu
fztLaZdI++IKfuKBAiA//qUEwnkEkAyQoQIUA9fSSeNQW6gAJu69wdEmXrkra5vQ
WGv1wLOYfyefVTl9PA4EFehw+QuyULSyvBhyZsgtfzs9vgaXrWZuilDi+dHb85SJ
nT3jOki4uR1KBRm1iY6F6MrtD34aBMifAg8kMwncNQKiVnyB7nzXdQ6PfKv0cZTJ
LeN1biOy6L9iuI2qyfzLW8tcslQxtq0tlIR4cbSFkcWpKNHSgacGQ9YIDufFpzI9
OfB6o3KfODVZVbhxw+iA/KlKuCqkN1ApOBSuQ/wyErFCbdkCwVPkKtNLrGB16W0h
/0TcJMDzNtHAfbMYi31AvMIc5q/CMgeJvhhP9FcEXerJktH99kPKkmMc3SAWxTun
4uF/D0Fs3Eulcq4V1ZsBpEJRsWxkjZI2zfYRhgB+BWSAeTRt/sxKF2buZI0ZcRIn
Mbwelon5jUq0yBWcCSE2raNMHS+2KAT2J/fuQN/AxHuTFoHPROnRiNrDxBLypqjW
NlaF2CHPaR8ce6yHKahAbz/le5PxBWVPp8AOovICuyp07v3Dgf/kNxKou1tLyeso
Nd49CrVHfZRJmVhWyPxWtU7HRKzCpsvo8okZyvWEej32gHVrEXxik2UvQugUGNcN
YtpSFI8qmNARXiMveL04S+iXSRPpnyzzHM8Slda2vraAyGT+2zF8FqUL1ugQ6Q72
KqQ7GZ0PHEJXvtD+HkVAPcVazv61sVdCACbet9OB97p4dIcJGclancWCpOGvRNHP
kHCQfQu/xfUApaAAu036Tnm2RHRWTeXcFczGHbW/7wpKXShk2knSEuGgQGGqa7d9
CU2bJajSlOWQTSz9RmNG5PIXuAer2M4yjgFLUAJybUEwFMvFf9nwoexUPKgdd5A0
YMUsT1VRKXweqRQIHXNsqV4o+1DUYlmpQ38jcnShCXryMkcbpS/svr2VZoe4HUQu
moFkp1rsxDqSdw3qJ2MKbml0PCIGBnwR1IeQ7X7YYWsL2en4pHGXTpqjQmh5Cyxq
DGeCwIHxQ2An3a91SL/7xjJ0mgOGYk7nzbJv+HqCHv3Be3o07NdKsPtfmaBRgJyt
zX9bH5rQqI0m4bHBWTfDxM5e1Jz29U/yqvdcKcND4dgV5OyPyfVQLDCa9BhBIpfG
fB+qi1Ktbygeb1vb+RK93X1wrQ7bf6R4do5rtFvNugdAxnYX3i90Ff5w4B3fOHvZ
Hk9V9pPB/HW4zLWlZeyeVy1R7NOMhHTsQEltTweW9qYnPRkiWWj/pFxPXxVHrMhY
eRoLFe3vE/CpngEpjEcOLyJae5QtWLW4ujfpdYSPjs9htNMUJiNii7U6A4KRN/8F
QFmj7IwgogN1LrXalVwsqQIIlTR2AgWOP19QA3KP1k7c79hGay9mrr9xX423pFuB
1On5mGiqIYqf7bKx+NrCSwy0nxvGeYHeyzKoDu3ouDzAZzBLUq7y5sy4PYXSsLET
pZOSWDV5VLjAEiODCsMP7D5lEkwb6ZP1nVHlQupS3OdkmT/bywrtfyCpOwaNVtSF
0OxSQynhTFMzqILIMhU131nMtcL8lhFdMN9Oog8eCZKGpI2hrNasecS8U5w0NVQY
AtLlU2+m4yt2/OmOVzYHzHwRRI7MFKgi6bFF0JuMc8Tm4igrcWUK8nu1s6vIbi5P
OuE7KFQB7QER+kp0zpQg3qzz34Wupa/fkTt8ZsVIBPvNwQlWXUXvv1SYrRKwIDCZ
ufPRGOiWd0jmTHIj1WVeZ0Fl/lg2jM0v+mjCr+1elo3JdbTzLoJNrgNgr+xejeld
Nxt1akOpD1pJt37HXizLK154sip/lJXnrMWZky+bTMskUItceSn5duwoR7t+Q57y
+A1aBpT7oJOCOk6mE8equktyT+6gWPjnOMLhuvnunEB5/kwBzN7JATTPX7qOnQhd
CjwtqQbzKEofc2MgFtyy7Hp0UgayJ1w4wsMattG7S5Mnhfvy8D0nvubXWXyYPvlx
zru853tp7zq65rNdENfN1iE+2MZ2ADOcuegO/O0ubZYjZROS9LPitAJt6R617CNW
XaH2GWUpTqWEnA4oacgGvCTf2RQ6bnpyR4yClWjEkO6vja7rQZHSjkrkQqripfRz
Et8rVQTwqPWGlsZocGViuw==
`protect END_PROTECTED
