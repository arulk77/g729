`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zUrO2M3R198nfKwSJIPU+8nka6vfB9uWAAlpUW8IT+W
9ZGpJl2Zdd4oeEP6pBHozMlpsVEr6luxSwp/fDhO0oXo2Ri8Nb2gbBFbvBWHNKss
GiCmZgAjE5hchYuW8k8c36AGnhEXKBuzE5mogEwC1DCmSoioWefmp/aOVt3yWE0g
abfaoEfUe1EEAsaUcXK9sWixJ8bVuIgKVG6u/XFGI7XXDd+tnwdUWWdkMpmlbkOt
a7lC4wPkWS3gkct92sbqn343UYRZicY8/KG9DtnU4FuHTIU6p6KA9vY08RJpVMYW
qse4DojIHeeiRIQqQoJhIby0cDhlu9piRqtZZgxq7/znjn6IjAQkpLHeuxRUUFQa
f0aaIbay4mHRit9s9Yrurq9yV+14CUlBazYYkB8vdUOJTx4mJZupb07r75j34ZFt
ht4OVC1gwqXJ/8yXiyP+YH3g5v1D2L+RQxfZMKX/rHyWWhhn0DnN5TnldkdqNLoM
cqAY+cUygz81Xkt/CBVXKflmvzEvN8jlqyvDv+S7OaY77yHRNlEK/dL9jG8Ixrp1
uRh0SIfqdhZN07vTsjS6CvugfFmv1mnKc7mZi6XMXswwQONbpwAUF+5JSJUAKK6H
/50xLuVy323OwrMPSiH0zuFhRcYSgLomGDnhom0DWpuJn3ZYmqfXNbNEh8EZopEX
5ZLnaxWrK8UBOpND2hZjDV9w/HsF+pRAPGEI34EFfHRZEqpX3oun40SfsLELzLBn
Yk3Y4lHp6NvlNpcWhsZS/f0rkG9LxCy8SQ2rMO7nZ4YRbPNfk6T9XgueQ/H4T1Uy
hBFP/tDwia5BlwDDyFw+0zfmjfQJq5dX3sBRx3KCxv4yL2dHuFMM/xc2zIC6dxLX
3ZPFvUTy75kr6QYieS54UTlJ1ZPUEimJfevfzoQ5gcW8XHaTTO+zV6eZ72SBXS36
ZPTisiLRTRmPSug/Kqf7U6IUijL70OciuwGLeNoedzewZuu8A92h1J00x4EVMKEb
xys5KrY+xVtcgWYaBgrJ8OztN81voMFIVcZoW4pQ4xWAwAA/d/e3wPUX+D1J+Fhz
x0l5YE0PO3RQ+IjLBZwvLWcOKRKetEbiCCqmPjjPiZTkmIaGCDbtoL6zzoNWsj5/
3FR1sZmsVeWy3TDGJ2Sehqzxr8W1TmQjE1LgquNOYp+5VtkzcTyO2bjNC9u0r6+P
v/8GkIdZqkY2Au+c27JiUfqQ07sBrAzmPxDTIs7ULbPhl1y0/6ckwpCsUFQ9J1NF
tA3pp/3dliRYH/H6pB5ie7jkOWJL2UzMB54oa3vYTSJSngoEoOxS48I1BvIaMvm+
X/IaaPv4y6j1mLg9n8ffaoHdQ49r1phDYp3wHZQlAVGyl7Dbw8whGJ8Oc1G7iUP6
IC3FiXHRMgK3K71F4BRszaVMShvVlpTIfpsH7L4zeQ1kx/sBsi7ciV0H/1bvDf8K
4rPuw5oa3RIqRzOTVAf+sVSWTsQoS8WGOh1JCrFjgDm6gHWre9hMCuGGHpkXZR9D
HIwpEtGb2XAMAOjLk4ysWlN28FLiaS0G9YwGbCKEJxCZuCjPBzY25zHQCXytNA/r
DDte8w3SFopUKrz5mrewB+FwuBXcrEA2VTx1WyVzecKVhUIVvrrrSk+Xy+B0doaB
B6jGQK1XmAiRL+u4aejcyHqcRo2+1jXEZokqqW8E09cVcX86mdd89/pbNQoof2V8
cmRQ57LL7zATnlh2TfPDlYoqaBPxTQGg3L//2PmnhVA05eDRuq6wUZNHDSoLOYN0
c7YhT8m4cUUC3rcEyAisGt4+tmlmK8MH7pyrXIJDArGv5vaGxPiMR/Ly/40cy79X
29Xhjc7f8C1DyI703iyUkZxFZdJNtVs+qnesIt+Kc4JhoDWAyXTZYnGiYF44IoCt
Gpaex9uSEbHPDuric3ebJLMHxwZQIItCCMWM/7O2o2waQY5blcrwnk4YAc1LQQwQ
j7FxKcN5/wgeellpY61LJXxne4j3AIgM8RRFZ0GsCpwZOSh15t9mJGD47Er4/OZV
Nn0HCf7uZCzIIUTQYpz81njHf6jPX1iMuNjjc/9WR8X4mpA2uK0acE2ML7Dw3eOB
V+HkXu+v9nR5vWjcid9tvYc2LrlNJ1OrBstU/pohmKTZbgoOtRSc5PnEKF1/KRbH
MiwqadRzvwRLoZxWO7+MBF/tTeOUcqMX53N9AcJ77L2iV1XEpPeDOjLOqA8/B8O2
r2/oXl+6rE8wB2eI0m4+Q1p4lZmvguSvUQzsvcnWFDw3unoADh4Zc7YF3CWcJQ0F
F0V7HuRT+HbQj68t+fE6vBWcIBZ8G3d5reBxsVZBg9dN3cKiQdns2l7B09cLs1Tn
rZX5ur0tsswAOvALHasmmHWhMjII11fUArSzZbF9JL19ol5MT09DHCgp2+xmvK44
TGN1u9Z9AxfjFddZCMdJjOIMEblSWXE2/sH7wyLkspkaPCRImoMFqcOYZy7k0u3w
rJKAokf2gQYoPKtupm4s5I8jCaa7oJS5XkTLdhfYKZ29PoY6OUREYpt6g1lOF6/r
AEMcP1H41VRf52HrbTCzR5BqhLJMlzCJaem9yvVP/U4KZNwHOcizgx4+mj/pyzLj
2GYGg9XdweXl7F5nJCYAmVoifmWaqaeaRu9E3oSYmE6jn4vKAsZM77HAzwULzdIz
nptDREFBwFPnJnJhLZn2KmE+cgCur/5Nha6lk0g1Jp6ajSKk2WHE2v+3up+PSwPH
Fp+IwDYlH2QdNPeXDKrFpibruUPLhyREoUi5Pe9YHPOeVO4mF5hkokgxfwsAzLE2
dmladJUYMESAyI4n0jt32A1V6OdKvBQyLagkh4QXfbMYcq2Zp9Qk3Xu5MsYAL67V
zaB5kp0yjTI0Nfc3KLSmfHCsuIekx+9Te+XNWp2nBnos0KHTSL6EYN7+9W0mdmwc
r5Km0ZfP/j8lTRiu1RzfnSdIPXLulrMr4cXpc6RoU/soRRc3r6mEeYgR35AxbEAK
GMSywT6vrrz3M6inMhUIJl+ohJY3MTOHVT6ZtKzPEy5Qe2WydBQVMy49W6ypWXRp
O7GdAeMDPvzWrau1UYSKBE2AbY/a0uQ7TG3Y7CcD/P0cPMe4zdrntKFcNhvCv/+u
wb44HFrt3QmRDn9d1CzS/JoRE/wqJElF3E8NWviJpuUrLAEnzhG/54kuehZ7LK5o
wHY6ryDr4m0NC1SAkObWRgkNp7Ucd5ePHYzUcEo3G07n953c7lS2DgHjEor0Ubyq
AVTogmHGNEar9M1DcdxCUJFTNjEewu4QwQblO8B4AyqDlbysPpOl5fPqMyLYh9lh
Y2gD0vZblZEylUog0HuYYg4U8M5Pba+Ss0b5zSfiw01L71l2YzaIfMA7jp1OPrKT
9WRcGMl/7Xlhci7rGkkgYGpy6onwNlUjTgq4Or74llmL/F+3dchohN/RAJ32nHRA
P7WkxX3awQwGDwPAmW3Lg2KRHbNP8UWsj/wIV064iYqRfbPXJ88zdA4E6ABq2xCa
6RDHy7NC/uMTiWeLMLBD71z8jgiVapNlj/ONXhwHPKXBYBxvMhQJ2ntqlB8J+2jK
ClM5DyygXKMv4jGoOmE2yCJDm6BRWaaZchvOOFd2PC3z8KqYYIRn8ODCbAlR4D6r
4atyxVidwtnoYtBq44MRogkRc2s4QStTHeLZj7nDiAz3R/VYvmed6s5U/YveLIUv
pebC8gLHbMyRxMsWJZkzLNTks+3xrCXT5Bjnze1IJwouiRHV4Eg0A6/T1sw7tucy
gV5A2TFzxjraVQHf7vTxUOr4Ic3xiKIHYmVMONPVn4oOyZuRSmHCiiNmSv67kfzE
G4NdYk1667PMxdm9DVeMv6ZcR9CHYlNd1fmbECGNI7p6p2zkXxaOQJgGSHbxbZGC
qwEVeRJptF2MLQow9mG6a1xNPLb1t/PQqAYNqzA+plDspH3PkjN3S3OaytinjFr7
7FA9jq9SAEq1DRmuzG6w/g879kQC5eVTqChILgpbUHo3uuQsrkTXVKPyAqEW9YKt
cV1VKop672mj0qiAlb8NmqFI1uI/q1lCZQEfOFIMEKOptGbN6hL9Ca4BgmrGthJ4
4+yL4rdMJUFm2Mr0wnkfTsTm+DVjNH9feXFF/siQeWQjjTTEiISo5qcszjWttOvD
MY5igli2BAM0gYK7v4y9ThMK+Mo+NAmG5xzXL4jSKwTzGLEzgA11bXl+D5C0neNF
ml3SpBBUnFRE5ljy2RmgLgUz/2RCaO0hOSNVfEjphbRhQDMR9PM1HxdbDj09sTaP
Tk2DDzyWIYKu4tNhDfenJ48f7AAKP69CjIqLjuea4X3qwJt+6Qzx7M21X3GTE2i+
1UG0RlpXn1x6t8Rtkktrv07QAG4RCgm3YeTtW6YObGK7lwbPCwrG3sqN6pUAdc4e
/WVvT+0WHtm4AZtBt9vivt9o1o9hLWj+V+9GB9i45yLytvknuyWAcK0mQ+U8c2A6
Q+rglDTxqMegVZ2PJU2utexUm0NERmuct98VbWxYMrIrDErG6MO87nG5vR5HX9o1
gRDtkzmCL3cwLzShbkZ3u+phrxIh11qOI10TOFPDEcSzbh+7Ovfr5UWM8lAEm3Yh
tbdo/FlEPMZ7HRkNLMBxReidm/VE9Nk8nKYj95r99OUzvImYQTZcimDAk+/yPce5
7iLL+Z7ImBLcqRM+Cgi+ECYK0hb+G5/KhJA+CHlraqqGSgr7x8vUuoRNsByaeiPD
jYQvMmPobi2DY+Sf9WCdlB8p2xh42IgfnxHwq8paG2ttGE6DMXdRxWQrbCDPGDFP
EGfWH9bcyCbbrEyNwK+LQlOsm3fmti8gHbL122XUf+vUDYieI11xDluRShSWnWOV
QlPxKWiosRaRhZAuZGkw1+AmpaDFsYN4Zbc6QkCoEbX80tkBYGCy4kvlFJ01OtEo
daliytif9KAxiAdSAyLRrl08I6413Xi4ziJw7plixGmluhG8hKeNtPjDC///vv15
31eYC1uf178lu4DqACfmca8pyud0KukBpuXRCx5BccHL9r/71UwT0GZZkiLaIjF7
JlHt47h7SKjCRjrKEv0UjTFKUupqbPHdXnrFxRb42vNV+3lc08Vy29l5yDj0pJWv
W+1stLFblUcx9O7sJ5cgOK62PJYXa0C64LfUyCL0/8Jf5JXmwzRI8qKBT92H3SHA
NoUeJhCjBd6QhysnjG9zvDGccjMxEd5kNlIOHgS+wTYQLeVwfBky3Yu4JCQMCsIx
X2InjESw8vAEp73Gb38IQxzEvLaDZ2Z5YQTXliCrNSAe7ZXDN5SGVv8SSi1q6ajg
DtCZ+C3PGo8nXCoWGb6CMtuILQ4/nIIZ4W3CNvgEhblfZxhhZ2PLsShK9QtgMIzd
vIbAwlii7jJ/0IONEIybvQLbmfVHbnSiCmzKLOKJUFJrAtJBSnioM1R6Gf/B35Pr
H875jtkCfeI75KLi1de/6kSzzIe1DR6UvjqKH9rH7G0I6jtwww8HidZb1Gj7u4cg
v6+ZsNFbM8p+oxQSEQxfD8nKZgr0wKm6dkKuF6LgzACuNLfkLHwzKWUypKGg9s58
TaLQ2/Vz/pXF0w8f+bWvRRdYu/6Cx4z857esjuQWxLNqjwKG54CgHEdVguOIYcBe
g+FeysbUKYE4gbASNysb4MFHsHiRswaziZRMvtUitzKLWssrC4+jLSMccyRmdby6
vRNkDn2I+rYQhOB9ZUT68JA3ixhFyongjw8KzXDH93roozPcttQ2iw6OZpZKp9YD
KO3G418NeHzOCcsRjkrMFxWGA0fUmxPwaYG7iOhMRJTrTsczH+L3US0jUj+FPRJI
esLz/QQNIt7yPtY9qcP+G/BVoTbLsC/Ohkoz1BmG5IKJlAgiyBVc4ennohw7D3yw
Smtb0N4YajaPqCqjYmIYAgCgc9wEjuE80tpSArDIxTI0gSDFAzWLyn+nVwFquZwG
bGouoNaDO5KmnfW+ePoTZBBS/fnRcDaaC2MfQZdXpGj/dAuLR2h+uYX+vXQLlcIQ
EYaY6uDnPGCiAFl6x0W5SJBUpoNWYH0yeDZrrr2Yl8ELP6MaBA++4UGVTFOQvWWA
ALzqoQ07WOQls4/F2A1Wx6jNr4+n+Z9NSCeSyEo6AQwPzd8JLUvgiIUO0gO+nk6Z
nxBxdbpWT8mfGyutBiAUlu2e0FYUWtosKgh5nf/d61mGoA0iMKb0peJBuIXr/4Kh
8UDVhF/Io+GTvjUIE+m72UxEOI7GT/69YNejM7u//PBt/WLG5Jc8WGVGZAkuVpp+
DElK+zQGAqiYEriobPR6RnNZeq+irJVG304eA3YjFE0LJi4gNPJQQI1ybdLrmFAo
+CXmtbzhq4nWKOXJ8fspnLQF5XmvFLK/rw6yW+oChYKfXhiF7DeipwGf14K727F8
du+G0GqthdcYsBORnswIPhFiPEkyo6/GF6YE6ujFGqbbStyFnIZKvuBLyDPHsUux
amExNhvk27wbU03aP2rBPPlD2yvMZzcPyPVAf6dqFBrBmvDae7abfC41Hi3wHcbE
EtRT1r7TvQAtyfulw+ObwiHHK5WfCVSC9hkIzu4fTBoY47NeFRyfF8Zt1/8Osj6b
cGRHLMc2H33v6dodiZSiurOIEur8heTP1/RfMMhGQk2JHz1h1xO1TNp1moZNwIq2
NhGPjMlWXNepBipfughJGvITMiANr1BsW9YJDNMzheNS2vsOednyWD+VQUFE4Nvc
cC8Epa6rO8C//76X+KDCXEN2osVY8f5MhDxw+Tclwh68NAl0A2x59BP/8IOhJvNp
M2SYe/smS5I0ZwsI+KJO6ws8HyNy2C8L6YvOgnLHkIQxVefQTAr0WuZwGJJcuOs0
QUf8Z4gF2RYlit3Xg7WHpj+VY9n0FZ24hL2OKQ8SrGhv6v2pLLIc5iPXeO6kUJZs
paT3e+3DXZVVKmeLFpd0/9z7/9LMQeEkZvQ2gd2KlQAC4E+WoIn18aui0AewNZ/m
LMSVSe5b2sbEEi8H/lrCmusr7sQGRopqGIPFfLaMOkNOTD3FY+Ltt691JpoRQ4VG
4VOb1kpvKE5jCDGXIDJbK8igT4NEJbigyUZvblR/Jp/zas6jlEVgv7z0z/Sm0AGq
zbd/kWNzXGXQKAVXxSiQqkckpBHotDAtkEPv5nvvY5/ALdTgcn3zNOjn0ueqek6N
`protect END_PROTECTED
