`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFdn9WEhyrHKB/x15GmEIv7DjcoZZ+3c+sl7ohGfrwVB
BVq4HU6mnblLV+HiMACqrjPDMLuPiFO6vAKqSt69Jpg2sMzLS11D9fu9yavzWwJI
KsZns6bBHw1XZQLQIcfzTqmUc+h3aObWkRgvkgXJXDbtr5X6Tk0EWJ2R0tiJ6aIV
WnG1OIg3tRZpA2noxy75TdMy955xV1b3Q3GmfTWaiNQPmadmKkXESQ6m+fqFl9Nn
x3oVGSfryy4+mAozxJR3ug==
`protect END_PROTECTED
