`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ai3z5HspTMrful8SjuhVkn1+RDgesfRzaq7a6yVdROjrYd1sZIj1NLmAsxcbXuBJ
L8tF6M1PkUmLodQhYI9Mz/Q0p/FNdzkxbbvu1I/jTWFeBcLKprE8yga7Xj1zo/uX
83w7UeWpEJRuFXKkgTv+z1QypXXq9zRvzDZSY2ITDQxPx5t5uQK2YgjQOcw+iUva
AdiFEsBWc5FlTISd02eWOcoBEcKUPcKoXKuwH9IJH2S8RWk85t5Mod6te6jzlb5W
diH8TtT3X10ItEdpwRUKVsN8C47gjZ6ppvWvXGq2b39zKlQr/jtXxWiVy7uELkjB
ENq4cOt9U+hfqCzn+koowCxxQyeLg4iL2YaXmEy8d00tkGZF4v1+XIlJh+K8JT3w
w33+YQ1nCdfHk5NXPESZKE83+N3smk9aGXBTD61SkVfz/PzLpVKZmINkDVcFO7EN
VNBCeCis5q3cO91Ab19QbSI5+xISj26Z8ot3sajaULaSJ6eeQ22iZ4m6fg75cg73
qsPyIV5HdJ16YYu9FN+RDm3k/8ae36rUhqHccrv2uiNDKufVVSkW4rKxFkGLDpp8
w8uKnnNpNzzzMwOPYCVgK1L077jCa+SUzzu+qVEuUfzBHHHsUkvzhhfRetbhO3ih
fJHyZ4K/yW5oycaAWOH24w==
`protect END_PROTECTED
