`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2TnjHhOxF+DAOEhybjr/y9asR7GK6zozQznRe0kFZ/bQN/M0GAT1ahPhwuHK6Tgu
fF5rNUeSEqWTDRp4NxBUOrEcaDRZ894+bOfarCXccSFCrB1AHrW1Y6VWCincJX9r
uBLzOWXJ+meYh0vIEkg90ShlohZZiOcDE6UZbPTkb3KLfkcR2xMLHUG5YIBpD2yS
pEF58+ZrLOUfDfWrWEWOlTxT3v7+VgIapvvy1KSponl58/wxNgWlOWByAbtLPkgi
CbbcSKP9S2RkPIswVRCOIOkb0dKKzwxxWWzUY+aGGqBNDavsPppP93I4UhYF2GKe
g7KD1Ritb32IhkiqBFn2SqOzqRNVwIJi6GvTo3M4/RBE9CxfEwpg8WbFg4pg32lK
UA2vobfEN8EKdmAnxyF2vb5xIQE8nY+0dnelanJRYBJCIRM5C8JRvznihB7oGFA4
XyI7V1fok452HwDUjLoAWA==
`protect END_PROTECTED
