`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIxlgnM+TF8aVK3WbbPsiJ0EnxVgFDnLU6d4JdTYnV2n
CX1iFdFb2BrT21AGW95Od4XLSYb5CKPa+nQwC4LIPahwZ+7oEX1RjE/0sf4ArlvA
F9AcDBon9kyNuYmXSc7HIAJ8/cCugeQ4E0BEjDjh15+59WPGQTZWOHPHGCmv5DyL
`protect END_PROTECTED
