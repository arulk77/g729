`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
gHbLw4KhCJFpgDRcVYgr8JtjJmgAH1hSSAj+Wq16Gx1W72Ee4l3mNRAfKkhWTm1h
zg9qNjlGq7HCqtx5lXWsHTQ7GqUcoGoiZh+FQzRciwNU1rUC042a6xDvBySTKIzb
humPqFFNJP2jhT+LuuhPGTP4F7XiU0X/zvOrtbqJyGjw8KTWIX74ZgHymNl6ST8o
ZGyJH37BDAeIkw1T5m54Z4e7mbwRHeBhixhV4HJbEWZYgm16nxHRcdVJsjSjq6jZ
DQILW9oJN1i8RXfwz4L2syBH1/johlngu6n6jayiP4xfaXkMi0IU8SDjuAoc46ex
cxAbJ/i2cpdv/PjfLRrHdLUqj+K9yDRe2yX5QUKkqRLEqFyId4HlxR45VZzc9567
OcZdEtYvd4P/cLi5NoOTtex2UGRhj0mS5BfhpmqZm2L9Nd2/+6vrYGnJAB88o7ti
++zu+8KzPwWHJntYGCSfgSHqYfptsFiUdWIUAkgXGpBlqb4fID1mXsna21c9qwVI
pm4pokRBaXo3vaFzzWXzzpw1rFD1Tp7kN5mIFOAEQapwRaxAfUYPV2fP3PIbaII4
eu8mcBYlbSjLMDFFyPjzE4V1NHCUs7wnqQif1BgL3T+fpqzdh+8TBoJLcBAqEJJB
XbcBXsXeQ+dsLKorxhiVgkn5r2Q4S2weeP/VNXuAiP/iNrsdzE4rCp0ZSXXGU/9V
0O7h33Az6x7kPbeC9Un6Mhq1VRm3zeQZhnLqOSxKJXcDb46NsbVCmGBikalP2mu5
mx5cG1ZA7DLsV/sL8HzLEmg8VreXfuURKpjx0Y1RHtSuEP6c83Q30JWDFP89WWUM
8SUrCWMETjN/A0dtROURl/K2WodFjmehtQ/85fE+A/7j/WpwK2WrnUWptt831u4r
abZ8xWIW6CsUvT+oB0mBj7d/JgmgagfUFsvZ69cX+qVGwWQNiMtFU01+bsOaSd+C
xqEJatG2Ig9ZJRPH4jCZZIudFk9vBa2vVX0Kp0FD16AeaEMcj39oCALKJsZiDb+N
jrAu3hOLlKz/Yu4Qz7pGocQB8RFJFebHf7TwSKt3TIEmFqCX7223QZ/2qcqZXY14
XZ7HGLkZS6OnWTf6NFSeShZN1NSdva1NrZrigLf03zcTrxwpVQAIWKv4Zj0y/r14
p+x/+FwUqWnJk1sLT+WOftoNE8M/tup0b7429RtKxJfZ2I8Qo+38T5Xb25fZEQ6Y
Ccfpt+WSzHP7b75p7q617g7SJ/0X/Oa0lypqLO3jybOU41LN0r2hBdzWOr7DO/Zj
ieTK315G3/W0BSy7x53sjXRWS0HoFlm5yUAS6S6Rxm1zxv4qCCkBTlgFvb+9df/P
VpZhMniFsDgYqOE0xn5Fm+RRz0h/VREiswXG88PHc/oe+XWwlfIrBEZeRMj5a+TW
9OND5zR1z+dwmwGNiI0o529pnjBpUVUoMGeJLAhio/OuupnLKQdfX10kPZ0aUaGA
JOLi3rLfJ6l5WUejze+XOHClROax0fF5VcnCgouZF556Hcn9iwVQ/cHmvfLEGhqb
Wx8uVqmEqBsWp6TMzDRYuBW9quASYBEm4O26g929Px8kTilxE92u47KA3uR5bDyf
`protect END_PROTECTED
