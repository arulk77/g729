`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JGqO4bas7G8YhiVzA4nkaz8tVqnwRYRnNpaXX+BbSLND+sgiF99Zv8t7ZA8KJOuH
jD0uGV0nkkJMV/b8Aw+W6dfyw9vkGHTBFAH43IsrFxv1Skkh9AtB1rTXtWOV1j2D
Da4YmdEcZQdEqrtx8qr65oQRnwbiHPeynI0zEW11xJwfIgLdPBwbE1Xn4g2LA20G
XeoR3H+rdh3/L2MQ4I/H2WxEVAfVOIEWutH10mibqS6O6s/q1qboJ9eDcKtu/ocr
crzL6ypXjAoF6rWLCmxZfEjEsAcPzYntMOIy3Bv0vJYq+AJUH+xNeaOAYL8EtEho
wDMOcsImfChAlYMFTdG9poaJy02Ehxf4807GKteUWjKo6ybwnSnaIrVGnfQIDMua
YxpBZs6vSL597gRIqTXGm/wL6JrkVrKGiEfDbQ3uYOx+fPxdNu2s1dc0Dy8Har06
wqVYCTCQ/h3zUAC2FMVxEfZi4v9vLMSUO2VOAdvMniexiOYVaXlMwfjuOuLd1QUQ
4ovbg5x+xrJIDS7Gipq5oHcJ8CQIJB/e6yFIO3Dco2OoyAu6edBpbDnzCKohumcp
sOh1s343PpZZD6AVrJEO4jUSrlDQOh0cDCe8d1T8plAosr2jZd2Yl0m4nN8GksZ4
UZgVAzjZRcMIh6QBs4sgEVTxpN6/jqWU/wT8JWZQ1PcEkbmLhODsXeonpXlZexJr
qTTCsswx2k1OPt2W4yvUtdj7qZ+evgn/LdsuMCvfhXc6F40Grioa2+I49MBXazt6
`protect END_PROTECTED
