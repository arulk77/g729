`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41wWADlDMrdCZb2Lxp9iV0Kq0QyPMAtHtcCBtiYl7qd1
ZEa+vpXpx0pc+/3o9wAnMbl7LeaxIEn07DCsCdcpBhqqfdgik0sUE75LXsqVazDF
AJGrh6+OnX91RArxaLL6dcopkOsXr+BtSWkoUE0I8Uj0cxsE7M1tA0zIgzO+Cbrb
NimVoU19tgojeLhERGeD6yqi4bBg9avwV3QtkMhi4Wk=
`protect END_PROTECTED
