`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLQoNRRlsC/3jWp0MA/u/A1l6BIqtWwUfVhZ3hwa2tqs
nF2ytMSLdb6qzh6xus0sXKUFqz1tqSjVl3D6vFxZcGOGwFNNpXdFzu2Vc+njoRcB
0w7S2IgF95+b23jIhmg5EolWMyqRX2wkP744MLuo6pAAeMCtVK772pVC1h8WGwQL
`protect END_PROTECTED
