`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SdqGLYzefwnCkldDbrkRt8pWS/PWpE6koKgQZ+2UC73k
7Ao1sOC/zZ4zlIubUFsiojL2iXdu623LraxLzlApj7UjRjUdKhhZOUHZs8BJHiq2
mPcAzJTUfaiwSos2LT2uGzv7EN/gJa8y2gPccbQ1i+32j47qRrU6drWMGCBXisCs
p8HUZIFIE6DVcJTBff9WsUeNLJFtQidrE3ufJg7EXAH79mhMTMqH6VIVUuv+0AFW
qngfCTYgQPM4yQC/NbFiRvPUF93Uil0TCOhLvAPkJwiiPeg2vEm7Jut1KyCmM+RO
`protect END_PROTECTED
