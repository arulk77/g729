`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM2llC4O4ZDwGeaU9n0LgjAfLOAq4bMF1oEFlzIs7n1V
PhBRXjLX+Nq/5EU+7L/nBbxZo0dqQKNfEoesF7Q46xWarbr1jXZTLlGpgz64PmBC
+c0XLGbS44RxeJ0m4QrnUq7quLNmp5FURn06TsRDKICirnGrwsT55541gygEeaNz
IRgdPQAxJwxGiQ8XSisgDQ==
`protect END_PROTECTED
