`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHfVI11ILivoguC7+j0E1LQr7792auwXzKrRURxjiRma
eBGAwpPXY+6jYRcCAyHS/o8QlxM36R1q3Bahao9g2POsohi4Ra4saWI+2Mix4oFq
N6Ax8l7nLuExrK57k4eZNGyqp195OppBGNWBsO7buPrdB4hCTi9s+190wDqoFD5H
Nfjk8cMU6iHz5rAyYJd6YYGVLr509gU4/75HsiIKEzUf3IJapNDJfOZn8K3WBHW7
x5fR8M30usOfxfGBrMP20cq/PwhXRVW9Iuk3gjPXp2EAzGi61/6E/gZvXsor052n
+ThxKneCCmY+J4TOrk5lSHKuYssm95An30TRvXz0tWSIG0/zICk/QYYI2uKuBJJV
a9AzPDeLeVT9nv7VoVDc+LIoPJZS4zT07K8Itw5SEeTIH32T+JtQEh4FbQmPcZFV
f47C2ipHYc1pKl57aMRGB19yClheN73arbG+xZ0JKmTEqUHfJVWE1ELN176IkQAM
DFpssQjqsqATvaEGtpOKJkWhcOn3P6foVxfdzu5P9V85GqcMnRKlUB1m/z/gXO7q
`protect END_PROTECTED
