`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu458aabCBUZ0DUXLJRMoeopc7k6T6ZChYPfCuQ9aZwFPk
XaWocuyqifE2kjtX6e1EbXZVpt7Ze30kbBA+mA6tCUq5eBvIchEocaNDMKmsBnvJ
4cNpbFjxh88MbwGzW5Z0Er4GDBN3f0OuxDoMqBlPXvx8y5hXFc/hc1WaDmxvTd34
giJvmQjLoEeTAmWIZ8FMPEWFoie8wciPK+BjMUWONM6J1nunXsL9g7LrjGydN4Op
P+bTzCgJL6a4kbSA9GXPZ7LL2T8YPAr2rMnKKErG4xdcPPPAyFpT8Skp3kRI+SPl
m2HSNDUOSCxy/TB2f0SMr4egO8ubH2EjVsk5cwi6ADlq0oC1MwIR0wOIuVgBIVdp
OXRlo3A5DzScB0BcuI7Cq9YANaOic30REhWsPbDktHitKDgKS4k5EW+COPlBsmfm
L7lvLvUx8agUhm26BeAXTg==
`protect END_PROTECTED
