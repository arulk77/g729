`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMFlmiOQL/IW4JYiJIMGbROUz4RUGvPges+uQFPYRMPe
AXYrUdwkAwuXa650GRhYPLUqS1+Ok9a3MSLVAasSiPyS7N6E/WS2hborMItos8ld
b3wemNBb1FJZXn1rE/R0Ory7UtMNfzX1+RI3P6TY/gemAwUbAAomze/y7Zd2i8EU
hyjtXkw/2wmLPOd3zqwFmw==
`protect END_PROTECTED
