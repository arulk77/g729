`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RcXNep9Z0sxKW1qy3l7p10GJL5+zmqfWKHp9Y60kUmMWLgSSiV1KtrnnR0kYXwxX
hptD4coX3hxTPgFjm2l4x7h2pMSc6Kn+f6KDwo9Z6JHMFrXksy/hyuYG9Apbc4HZ
FAol2OIXGFnNQNYVkCdMG3SNxm6r7vI3qv/ha7nuL3rq9o8htRM3jqEIoNhNnAjQ
9g/ASwbNkWJtMA+4SpL5TIem0762rL9vebKN1s7+CdA=
`protect END_PROTECTED
