`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49cC2bd2gjeBjmpIDrs3Vmxj+PnYgrfGNcQPDHuQy0mo
NbkxlB4MzF7r2GF4XYaXjLgnNtRhKTGA8SVi8IFDnF1NupHykJs2hFxcHqs1s8l4
Q2OdZER9Dy7esNziopG1WemG9mn/N6ngC7E/Jy0bRsy9M7iNi/m+Y8325qxwvnKD
JccM8BwGdlQms/b/AHuAqY08NgIJglzYEzvIjiv1AgLG03uwjJHr19N7GXT8KXYs
dW8UHAQipkvtUqbMLysEiKXXwBERlIAG6Za4L+KCXSc=
`protect END_PROTECTED
