`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xJV4QGKNE/TmZ6FVbw4ADOACB07qNm8Tp2gHatJRgUh
uLDHEZjypO9AYcRh6zJFgxxoi15rfmmVNFzDFBThqYW8C7vxospbaNagofFQM8pp
Kic5QR+wCY0l297qM1qMOKLUgRzAu3RZ3sQiPGJdh2HGDgTQpgCPvu2oRKP9mKdX
+Fn9R58Mr8PQfnpwvZhb0r0Xh9IlpxoptHq0g1Bd5ibKIb2yCYvqr0blwEVajsut
KHlpdpFZni8OTbPtLCW4y8Z7a2i91AVNJk1Y1PzSHRMnBIYBtnMWtACCDxEZtPTC
rHiVZiMuhneHSPxhAK0jiZNqvGuvAsFgUfaNt5XbGCmRsh1tI3pnyZYvOdDj7buq
zvELDBkbyb8Mlg603nB6qKT30/0sO98Yr6bnkCydV1jNk2JSuwvpw0kZlZ5NKBX+
TLaQzhpTRK7ZfLlVJslxZQ==
`protect END_PROTECTED
