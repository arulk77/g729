library verilog;
use verilog.vl_types.all;
entity C_ACCUM_V7_0 is
    generic(
        C_ADD_MODE      : integer := 0;
        C_AINIT_VAL     : string  := "0000000000000000";
        C_BYPASS_ENABLE : integer := 1;
        C_BYPASS_LOW    : integer := 0;
        C_B_CONSTANT    : integer := 0;
        C_B_TYPE        : integer := 1;
        C_B_VALUE       : string  := "0000000000000000";
        C_B_WIDTH       : integer := 16;
        C_ENABLE_RLOCS  : integer := 1;
        C_HAS_ACLR      : integer := 0;
        C_HAS_ADD       : integer := 0;
        C_HAS_AINIT     : integer := 0;
        C_HAS_ASET      : integer := 0;
        C_HAS_BYPASS    : integer := 0;
        C_HAS_BYPASS_WITH_CIN: integer := 0;
        C_HAS_B_IN      : integer := 0;
        C_HAS_B_OUT     : integer := 0;
        C_HAS_B_SIGNED  : integer := 0;
        C_HAS_CE        : integer := 0;
        C_HAS_C_IN      : integer := 1;
        C_HAS_C_OUT     : integer := 0;
        C_HAS_OVFL      : integer := 0;
        C_HAS_Q_B_OUT   : integer := 0;
        C_HAS_Q_C_OUT   : integer := 0;
        C_HAS_Q_OVFL    : integer := 0;
        C_HAS_S         : integer := 0;
        C_HAS_SCLR      : integer := 0;
        C_HAS_SINIT     : integer := 0;
        C_HAS_SSET      : integer := 0;
        C_HIGH_BIT      : integer := 15;
        C_LOW_BIT       : integer := 0;
        C_OUT_WIDTH     : integer := 16;
        C_PIPE_STAGES   : integer := 0;
        C_SATURATE      : integer := 0;
        C_SCALE         : integer := 0;
        C_SINIT_VAL     : string  := "0000000000000000";
        C_SYNC_ENABLE   : integer := 0;
        C_SYNC_PRIORITY : integer := 1
    );
    port(
        B               : in     vl_logic_vector;
        CLK             : in     vl_logic;
        ADD             : in     vl_logic;
        C_IN            : in     vl_logic;
        B_IN            : in     vl_logic;
        CE              : in     vl_logic;
        BYPASS          : in     vl_logic;
        ACLR            : in     vl_logic;
        ASET            : in     vl_logic;
        AINIT           : in     vl_logic;
        SCLR            : in     vl_logic;
        SSET            : in     vl_logic;
        SINIT           : in     vl_logic;
        B_SIGNED        : in     vl_logic;
        OVFL            : out    vl_logic;
        C_OUT           : out    vl_logic;
        B_OUT           : out    vl_logic;
        Q_OVFL          : out    vl_logic;
        Q_C_OUT         : out    vl_logic;
        Q_B_OUT         : out    vl_logic;
        S               : out    vl_logic_vector;
        Q               : out    vl_logic_vector
    );
end C_ACCUM_V7_0;
