`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB03S60OpZ/4gGz5K4fX3i9tSe75kFBJwYBPCpTYz1/J
XW0m6cqOXl+NFbZJ+VkjR34leW1Pq4XvRs6zOXo/85Ye69GguizR5LyH7KWFtXv5
6y4qjdfM6c0V/tO5xptAlwwwgFiC3BAV1nWitgFgtw7vW2cn2Znb0uXcrVubZqsX
BNjPzm6mcB4r7mvQmlmf0/nr6YXCpyN4ErwaDWP+gKwsbsDGClogwg4xG/cl+2Pk
krgIJHX5KrBiG0s2VIgARasgkapIw4t9FfCBgAxtBg9Mush3+xPcRkVTjm9xhiK0
MmRvv9kPqt8fymLp+F9iCg==
`protect END_PROTECTED
