`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAXnNRHzxhjYAW+hlPZOoqloo/rwX0VYeMpY8Tx9ptDIb
+Q/dU6XiPTP5IpOleFA+AKqFLJ6Et8jmmPz0RFu9mtgLbQePIxdjCSC2OrEfCBrg
lg6XZULQeWcMnEMGfyemiJ6Rrpd7QBaGC/4DS0zqG/NhRXTVIZ1VEXE4k7J5xyqW
rDg6V6hnzcuWDxnq3xh91Y+dNW/InJnzwTFzxag4IAdEhuhbq75GbXg5vsYAa/ah
BCmCEYngvvPRrK+yepVXkhd5QJ9+uiZo4T5KRoV8nqqbnwIAnYxpiejabarOoljR
pfKyRkvXklkRJbjc56DniaFgKd0oDn1PFyme/xHfee0ow56rYCXi5SNygioWNbce
ro5E4NqUUdQMoXGCbsfqMvHMMiMd3xddZ//xUeHDe7hQ8OJxrgOg+SlxX0xjylWk
U/QJ9rY+/YE1tlYH9Xm8amtcUWZ1OwzYGsnhM5VMES0QrxsQIpCHmJL/DuAcNwpZ
hUiVJ47gBD17hH4tTeAqaAb9SFyYidCqfzIewvd99f/mvinIKt0DjG54w2zkfQuN
w327LI3Z4LYXfOyPrGdpAtbsWwk+ZlVtcE1wkzAyHiDZ+j5vTDF8OOQz/rdGVOYu
cu2carJEBOCx4Fq91eUlmCtn9DFw4FpoKK/wPSaZCMs52dQbyEImJRHO27rgXBt0
YmuO0o5sjjb29vROMuXsu9MO/9wAQobM+kAxhVqixWX+xhJBk3kscPAKIQB4Nz3q
sUrTRyp2QYqLxPjnbqsF7sUq+uZgDJlaiHIuSFydjKrQYaoFTu/+U7CRdi0xwQf5
PRcpNDfqnUDkqBy9pjjzCYWtXw3fve+p8iLRgXj6NDum80XgLvm2pWPx5zmu4lKk
xWX0BLndav+VXd8hxdwigpDRppP7nsMJTY58V6xE5y0e/SnTDDaLbp+pKi/+FPjD
pxDZDxkUczrtIx03I3UGKzb/I4PVhk2UihOYIeHHa/I63sawjs04vfB5UJOXP4Es
kZO9GjWnUEJr8O8JX/+pWnHiZWGpM/yKV20UrncncyfT9ubm8J9SQP17phN/WJHN
nDtyNTcCiphG7CUKdYw2ROs57gHi3v/Ovh5B4lQezruWTEUluuDDeFhY7bHLQPjq
jNDiNZ2uuteq134ykpB0vQ34uEZ0DyDmW8UEEm2xa8ZQ2Fo9COwOcS8SHoFKge5j
vkYTahoCPf6jWvjBVCvB1FiK9Sg8g+SCRly5BX/v3lP2TAZflxchRIiyRGVda3oZ
NOWq10Ex4iP1XWnlhZR/NnMzly11MhURzV9uqJ1RIr8WzefdkaJjNZPAR+UfyvVK
SWksNGxihXGBH5G2T6oMos6BSXZhr0oDWB3TriCnSx7DjEoHcuVbXEGlWt+JjWrx
U9U9MLhG7Z1UrAdEasaDHBqgKE97zaAFuDf0+y3LFulCUZfJbgvaT2taTst90Ll9
8ez5GBw1crShRBn6IJ4LHHZNGrd0lBoqRsHXgUyY55mchZTM1Ii8vVl8vTLRRz/A
ddMBFA6O/ByZlmJSSNf7/dkKc9TyqKP2cWYbzCtNWiOKv8gKgHgYEI6KPZqZgW23
IIyyyCpHd2LGimF/MmVHUcUi6/qWC23R/YOZ063GnuT2vkwb99imphUQzM2hWVx0
fvbkxHfORV496fbYsHm4RPOjD0+y1djrOESePKumQM4=
`protect END_PROTECTED
