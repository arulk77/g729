`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBbw2kdjAoXLXZcd4cnLfT+VvwvuJfC2C0zSqDi8RV3k
R34W13Aur926A2HHCzPBCeH+ccOgRZZdfy00PhHnYnfR/lqVglrErmLMpqETOeYd
Ab/TS9nGwBNN03NFYNVnpyo+gCMQx5xP5mim9Xx0PycnMqA8y0WfLYAKC5dyxOyo
SxyCq3dcKpw66k1L/kpROoRKJdnXdo8F80y4z9gSyJJq44MidKng/zwqus2iTR+q
72ryfFsZJeBr9GUtgoqFrjvI6TC48vtUcXQPqHB2vNp+fBmIvJcgS9krPZBAPr4D
j8csM04skIV7nuYOz2w377B6FQJis2sU1ucIDc49oI5HrAXamVSNgt+uaj7IvJ8b
DqKo3UEqX/eM38FPn6UKPbYX96mMwB46MGwVJwvxEf6kgj6Wibz9f/joEKYe2/gZ
oN32B+GmFImrXpFogzyir+K1rlgafZ4ID/o8cfP7v4sI+TgVVpgHVLNwM7duimP8
s9J7bTRdFZOaxmro1l9kEIB1V+cdGkP8vkSiFPsVGa8U0sB2nipf0ZVj0ZBf+QMQ
`protect END_PROTECTED
