`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXA21rgiuEO5yN2AjcKeGYKALXEJrPffIMr+B4UMCqKk
XzDYhIO0DZYCzRcvlilD3ZpmzlEl294COfg5kWPpdwJuJpEopM9BzO5YVXZuwmfD
uK/BJGDxN+VISXb9FnPKFi3902AhbNw8skDIe01bE3eSnKJi/jvHrpglUDfgcgSx
oxBrFBCHTkuKexETuE/+n+yCD1miAEFW1RtacabqRJI220OPbD/8vsksbr8Rih4x
5mRODFnxG08haQC8NziwSDETSbcEJzJ8eLWXm24Hg8LLnuAczN9jIgkTcwK3Tt6k
zZfiJRhwe37lAetU/KjL6Vg1Ra8UYcu91YSjjzewT88=
`protect END_PROTECTED
