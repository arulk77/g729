`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD8DDW1CGRVR3hU6QAp2hSJ7myxTfneciD1/PL/3qWfU
zfX1RokhuifkIdG+d0Pe6gDbLTT3qpyjfsyxHpJNTHiB3QeiqU6OdBHugusFuy7A
PB4Dyu/VHpxuEi5kAWpr1zfFZf5QqZh0XSvKwUwCJVNDGwF7LhDI/QLQSSx7sDsw
`protect END_PROTECTED
