`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKdzjYa2Dycj0cosOmI8CYimvvWqMYnxF1g/gWej4Cew
U2nkHlgbGtlRw+6W6iYX1cTCmvp0EvxMBtSJBRTJm71uBeyFTKBeFpl469gtFWXx
uF9rvqEVpdmI8z8IqfpVODfPgXHLhwG1+JRNHoqr3HsJv2go0p3xS1Rjl1KX/iV3
JQ2yHnsXi4kJn28HiXJA5Mbm8Duow6X8oSUkoe9cFCw31mtOvOj3jK/4M65w7jlr
o/kyVxVqrzQONIwNm8vWV7fWD2DeCGWn/gjO88uFWn/84wn9OKFoQjyBoVsWfnjw
ofUKvP9IxTJGss3dIVh09R+Pk2UqBMY3/jFpUUrft4f7aWhzCUSqOj4tzvt/VKyf
L0d2j+IUhjqmQTiLi87GShP+FJWfMMVEtnFGbXYK2pZ9LxHE8PEZa/YemIA+tv3e
vKAWjVO4HKjM+ahLPDc0hvHJc+gichV6nuffF1MaDXULOYmGXyG7UPs/WQNfKY0v
irvE/ye5gdTCm0VRDAC2H2ksRtr9bq4PHNVT89BQqcHlG0cNEPmO2qOfs+0Vfm73
ujbbW5SwpcZpQolScrV2R8SffE2zIZlrdoDl2rEoIxjI4uq5gUcvzP3sKlwN1Hzf
`protect END_PROTECTED
