`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBE/I+iZCDM5JuLbmOSb/1ANXUQKQgArtyhtXd5oH3CM
A+nH8nQjXcSRPZmD1mjC7xKi0Ff4jS5zKBV8RNrQ1RwsHGOSFr2bQ7EQVtti5lmN
S/rr647rhNpDVFhE6XoDaQHnWg9cN2gr9SUPCPdX/aGPSeoJWgpg+5X8aDrcAQLN
xlPDwZlta4vdoc6zvAFypgNGGBIW/ZOaanZienwWuDMnpA6BzUcPzSrfI0Ca73Nx
OEioUX11hYKLjTKKNP78TQhs5VH6NjxpefBaqcF2tM5VdTRGzgCU11Jqv7a2NxXE
CObPCH0rKz2pSwfzDtQ1zl0/JcbY+9L4pgSn5HqbX+QDubOMJykPotBzkS93Kk/t
Y1LUXQ1BylgBH1GaKozO06+//t2GlaEKe3J9mPjq5w8esNUx6/dSct6cQI0Ek+Cm
+a7MOrux3YrUioyRY2cDw5ixi/EfVZDng0ZCJ7L2/HKFNqAa4rwBndBiHitsa5CV
kFg9EC16cd6MDOhHyqqLp1GhvCdElKTpWmwGy5BDqtyTHXL8r04nZp0LCzydNS4D
gPoGJg2w1pvFmGhN932dp99avL196fxNZEPrBHWZMcETuTzgzERZidGP0k1FeqWE
I2eZlvfrJ45TNj/+AQYdisCr1HceStp01bXnLUAaV5Djn8P663u886moIoMJmXGo
vdDHerpBxQOuCYH0DopZIPndaDgnwuCTYl4SUMvlx7B+Ovhe61M2p4e40ymFckOt
55eP5jCgxSPU6STovmMyAXATvjk23HT23J0KTQ+Vsswii4olmG+86Zfx/Kq5rRx/
oMHZzAxy+JxAZ8O4jYecpt+63425ZZ3N3txOu5Cid9k=
`protect END_PROTECTED
