`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBXg0I5qluZrzEQ5pwiXw8hjHhESUv/EWP9wJo8azMnc
6QGbaJXdTJX2zYcucmOQKSh+Ehq3YtJHHBhAEnIsgqcolwj0opesa5KIImcNiGnu
Yfq0UMEaMKsRq7xOyd1yNurVvlnPIZvmbDKxTNUHgJgQJ5zLFslDaMr6Mt/Z/h1S
`protect END_PROTECTED
