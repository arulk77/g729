`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44n8kSTmRyFAb7oZP0G6PiMOvEJbpq4KxzHI1w9PU8Iu
lNysASDtblc3+DpfwfZjDvNt/gszzlC+Oq1sfYatpO81eoe6U992eThyTvC0ETkK
U96e4+xgFhmlhyGV3W+V9koBXB5QKfcEhp3YRLBszptEvt8UuoGzE3E3p9rpOF+i
xfxfF5/Sr17JiTibLB8p6/LitOwidoFdHjHjUS5DYf4S6x/4uhz3JjjRLM+yw/9o
9S9ef5n0Y+uAxxYZouo//2aOEKAJ3JHfyzPoSQWjISysOG24O661VRKbQ0FzWFrJ
8HYyZJWK5CZcHD+DgxK7ah6g364O6CsN0sdAPwHa6ca6JmmMGyplUCtUzcsDJxiT
MbCDpDbycWsEmIMNh5lBbe9BFpk9TZtMjA+U2rwxmdl0gjMEnOqnEaaIBRKbiTMv
0P4OlX/2BWrDkoZ+hLdySv37f/Ena40avdDfgZpY5G+93GG7nWmhJjtzeo81gYGU
`protect END_PROTECTED
