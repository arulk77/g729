`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKTodPHHVTK/6A1CKhtsW0a7y9876n78EVXuAYRm09Bn
uR9A4kMgABWpVwU9kLrjcWY9+5Sgu/8OxJYTitIV8pzXvlZEGm2vVAqYXgi+lHiz
BMkMUlYX7TaBOZhAeqDi7/nsLAXnPAr+AIrl3q2JaKdJdTWD94HrjUytf888ogXj
`protect END_PROTECTED
