`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDw2A+AhZc5/Cvty90e8qYEX1Vr+XnN0e/k3DSBP7hvf
bAF/htShyPlim3gKBNW3DmVCo58NgT9YxvWBp+Q9pbLVEAQPZWAQ+bGgmGuilW95
Suy3i6RyBeLlppo3nkjfScGYkBa/bidTMdH2AupHr6YdVTk62Lz4tOhHYUmgo2Av
9YRMD7DvpRrPiGS+YB1CApDMB5CI3VgdkbeETNy0O+xTzp6qhmzFsfNVBHKgIJuD
/euS8FkboX8Dm0hJgRi8bQ==
`protect END_PROTECTED
