`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH94/hSKTLSl+8CH8PcDJ26yCCSoOM9RjqvgwapYq9nL
Wbw+dN9KuQkKT2Lb6bUasFfxvmJC1AR6unVuxPNft7Avdfr4sGiyFHCe23YcFSXK
THmsLQv5Ia3FJjH+UdxCees9Iir5Pr3Z/UfdeJxux8uF3uJ9hjYCPH0Y+C5XMF6L
hvhL5FikwD4/CUvVOZfQVBlfTU9B2ZcwuB+3k0KLgDlmEO26We+1JdY8j74ifoUw
x2YrBQWmGumkFHxs3lTRj97EteFPSd8HR9SwomJrdBttRvnuFExyNN4ZGGEcAJO7
BgSAHR5AFzzXb+oC5PNvYDQExvKSkBqGv+oaceXgzYF/99mvli6Hq53Se3ZCAkKS
0h+W8Fo2pt7fs1O9AyfQIFQPO2dXusn8+xDkQC6FN7ngR7pwOkeWi+m0FzgiJRul
Gyb+d3ItRlqdCMM2m/omxh/77wU1Kz70rCxiYC8n8GN+jwKhiW7+hIxlcvTY89Qz
yvEMJvDaXMd+weiuqmlNOZOw0yV0br69OUV+H8nfNWt71rFrrKqhD5n7JphOYlFs
`protect END_PROTECTED
