`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CycXZseRWWlU/Rl8zR7BBcMHeKhc/Uyzki3je9bTOGnI
baiZbz8IOOiU4iXk/fw0nGQ1uqnyGGg/Z0AQCu92Cwsc5N5Nl7QM10MEf2W8jlyE
fjSTIEZJwYzGuVXPC8DQTcMQ76ZHAJJgbGNAWuL7B+2rzop9NXQeXhvxAKWHqP2W
i7VK0kiDvEcUeKBYq6Ib/da+41hQxboHWrSKv/Jb9VpyCJbMqdpn9txay3FHAJe/
yBVh3MmekR9JkO2lj4jbM/pE1ooMomiNUgzpCHPLn2tVmamFnbcq9n1ypCZ0JAVL
Vs+t4IiczwnULfPWT8rnVYetlv+nRZQ89xbPPs0kPuVg/UMJiF+jO/DWLBt77pZB
XlGbQfcdHS7UCzZRSK/whaxiH8RwOUgfOOYsPbd9oofZjtuUSXOcPD4iD7EzotgN
YIV9WEN25tg3L4N66pnxh4ZK2nX35TLXbeTKYmMAWfxq4+5BTcflyxSxdNLi4dIl
EgC4ZnQ82lNHKQx2t6kvMCj2fNCrq4RrF6kX4l5tDZIAUPW3LbHlcKrZZClfYZYy
Nac/OsMB+2eHYxVttitHrvBPrXfykKqV9dFBFS+0cCYpFjuI2NkQ1gkC12RdVeY+
nXNWU2TAcU9mvumtmvGFyGsplNA0Trrbm0VHXadnVc4zkzc+FKg72YmjOP16dm7e
NwqwQ4hx8G50HWX5eFyLPsS3TP+WgLVjDVSg1jr2nRSkG0F/eiDoq1v3B7gc0GT8
VnIFEfgcyecy3e0FAst5aQI+lhWH8IK+KyZ7Pq1naEf6S/mA46d8pU03MfjYM0HT
lhwTTzx+gwNb5IoU0Y6fQJlIA83N926b/x0gIUWlyOK0p9G0NyyEzhyuelyVS1hw
TXHwEgexACK0Z9vrcuqjGc+3WccJqiXWKiKKeXSfza0oaPJQ/QjQl0Ijf4gKMM7j
dy70Z3d3aRl9u9i9F/IgXi1rENbZo6I0t4qL+TFIcdykaxUOVenNobWu0y46UE2H
IS3YX4laVy+THmzc0wTJKcDLkAdctqtJsVYMaJWJTO5UVHKtoO+302o2er3lqMFn
6LFT3EYBnF1rNisGeBmr48QdxDpBKWZtK8y46ziOYo4Lq7GLyRijr4r9PHw1ZiiH
lXp/09FLAGCNCIXZy8H/Iq+RmVFb+I+9JKsGo1C2ltkQTL2xpodzkqxwc/IkuoNd
wc42jTcuUIgN9axFZIbJxltwk5lbL0vwzK2ZQMNaGEZLpkHgpeBP81ThcoVR61ZB
zL7S5LP/5gF5P/BSnvLURx8JY/ZRaUd4ck6XwF/u90fnljtPiq7ULDR6uiwyKoYB
adteuQnSuPpsOu32iyGy0qAAAsVFwNYd0BvMux3E6V2nZTp3EnRAAebzE+jcw2MG
pJatvQWBpOsZ3OOktfdwInU2cbZvDOq18SX1I/jD/WVFmm6m1C2bmSKwpjtG+vHl
P+msWCbnVvq4BfrYrQeFTP+YV5PqgxEWJewkyzt6dU2W4rjNsd732ifsThU7Td0z
w3sr/2EalAyrxlpXXihKxGp5QuZOZTx+YM3Y9c3VjFdg/n+GOWjWNZiVcT9P+ZUv
doW6SqRqMDLoxOJaUOhrUS6sQJ9kiz0qE5pR7zYgAzcPigrDitEE/kcOUqoDl8sS
TF962weV3QDZnaVyNfwyIMnag6/H2vXM1fqh/K7h/2HNJ+wHVlapjVRtZ4WKKmzC
3fpotvCY3K/gQ3W5RbeE8PNQZJyVUKDnBSLCwlP1Fng5+NEEnvlhv5LqID1rEnKe
JtCvGertNdy7OkN3Yv8Oi/L9TU38MDVIj1I6+ggm9XGpl4ab8BoGPscKnYwi1aO7
M2pLr8yWI19YLMCRql6lJYpH9XzB5+gsOr0ZAQWj0GVcJiB5oxhOl27al6BvR9LN
OerjCCMODy4POwu+kkz8whiqH2bwH7Hc86IQ3hibjoG2zfqUkYA82/dDFFI6PXBQ
KkfvSeqZsgS0u0j8lTN2fcEUWG4rz0IszELDuBbN1Awy7sbdqEGect9w4qD1qrc1
qBQbiiglC2Bc0D98BpjGgwSDWKuWqmigtC7F83bspGaE1Uzy3HC5FBahiAbP1lIT
tRqeBO3bT7wjlLic/sgjlFPl+2SemBMFAaIpkUWqpvNhlVyfQHA2ctWTZNNJlkWg
VuILdfPHTK2eYqLLpi0sQLlg2ZaZ6JgafhdkF1Do8B8wrZ9PJ7J2K0f9+p9NBf5q
o96yHapUVEnh4uijzu6wFpnguZ9skMv5kpi6+ZUxvvyBPYEfsDBjye4433lc4u+x
4mLBu0BQvVkJApYum5FEn4KsxJ8r1NaILUCCXTGJjk9LNGZieLx+jr+3AFQDI22T
cde7RX2bcmYn6gvUz8OgjdIJ89FQfNJhBfwGPAjLpPgJWzxRinFcK6/vBAreAr9z
TbM/UxpQn58csahv39j7z1S6GECaRygkdJMiBLAGJVcc9ouQOGlcqcb2kM5dyGY2
rduIbotl2r58Xr35W65jCZ9pR3Cg857qt7J1PBWzfJ8+ZurAJvY7Q/hYQyPt9+MZ
1AyH/Ku9KJ/hlnYnSiBA2JIfFH+Ox+otXL10NCvklQtOtNT/AdeZ47Vb0/iFoteB
TFrcczQy7Sf0eAv9QIXnHara2t/dW6qtkh8POAF/b687jiZ6+PC7et9yR5CGQwD0
v0n/J40ayR+xbc3be2pA/Nlb9cin4l6seMv2nKNwEK49XHMCN/ZXYbofpNRGRfbW
BTdR9+HbYjTDltKm5IoOl3eBvK/jtNsjdALlkza3J5wMs1ML+hQWTr44q+Czs4Xs
lyc4FtMVfQwsZdc3jIosRAKdz85krJiVSWzQMmbIPKXN9KbSnF1FET7wxJQJ53yQ
eRqAe8pw3u+Rtg0xQPF+/IqKX41+t0yU/vTAnpq/m5Ieeu5YCVDcoKv1GsvVkOrW
XJ/yoLuN/vHM0+7ghgCEjwYtf/2KL62KbJkcXEoN4sJvv+h4KLA19F6jkI3JHpFR
uGLiN7cPRWGty0uySD3350d0H81bYpwboyVQrCcJNYFWXMt0ViA3yfGONE6e2JxQ
UYTlKLkZ3jK8klF7mGg8fZJfJAOpc45B5p3H23DkWD4sCVK6a42adIMUIXhYwNmz
Pj7sbeC348KTd+ABuGjG5KNwkfejV7twjORhnZMFCWTgSTi92rVntWjeVdg7mY1u
drps0eOPcA49Twq2l2N0XbWMxwJIxyxvq01M+R0/353m+UMp/6zU5pndzJQIX8/X
Y4A6EJladLYW+4qhjZhqZpASN0u1bmh594HJu49tB3lXamZEDDsRHbOOMlAky+Ni
uBAZLudYI23mJSPsW2fr6nCbrdUs9tQ1wZ7qDHBbvE4qjiKyP7rI6iyenz7i6Yod
6yutqhz4XLgOMEEmXjybucoxqsWIa6I9xlst9mX0Ka/2zfaIh8m5L/y0mbkQkRjg
YC49uQQygfBeXjbPHRAEWrR7H36u8HxM7RzzKH/hjXZsVCj1IotjYRTIpsmvVeyK
OrCIvkbbscQn0LhXAz+h4A9r0CGh9/CNIN956YLX+j4e8Dp3Vu3wuLA09Ev231Ih
hRcPWBStnx0m8NYyK5o/7MKquxr+/K9/KziVca1Ndtox2UOxpln+ILngOsDq4nJ3
I1tHVQCbu5lgzC9PKXmsX2wt1SuS/+i70T1wxH+Y65N6d7tmCEGg2v/RftMEZfIF
`protect END_PROTECTED
