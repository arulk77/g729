`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveChl1uOKRyac6/g1Ag/2+S3JcG6/teKLFjsxQdV3La9G
CF8H4TceR+pa4io5SpwtYrrDX3Y8WSMxTFqdoZBPkb78vfLx8MaZmM5qjaCRqXIy
E0Dhy51d2V5dsF2jCRU9vx4Zr255XZIaLtNSujGRWlyQs651pB1CLdA+GeAhUV8M
beWTOgfJ1Wo7KR9fvzm85vJdUCCjTav8kJe83NNw/0lAwhNsxivzVCDmDw5c/ILF
LxMxunettewIjQjUaqi58SA61hZYAI4mpVoWdkmbjeW0iBNIhtzMxyInXVlAXE+/
oljUQ6v2bgD4LLj0cROBdiGtD32nDMmpybCKvtDiYPjcGdFP8yVQq47bjdd4/UCQ
oqvpNDxGuAKrI0T3BAndRA==
`protect END_PROTECTED
