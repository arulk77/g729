`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GiBTxzHwh5QDbzjhnYEo+gishv61Lq1AKwFU3oitGdTrSv7KyHUhC6zHPrecMars
LXxwooghLSaqktCAJv+5B6LbIi/0wH+Q+1oWnl7xSNH1RYHJDj0LWoZWdPrWMlo9
BXLLQhSN0JbdLXob8Rk0IeLTkwyW+A17olZbhv2/FoSrPU/2LsOrTZhRUzjOpF4M
`protect END_PROTECTED
