`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePo+c8AmaHpqmblhcuismYxFzUvZcx4KEY7BX4wEz8Ek
TkBY8boUkffkkdimTUQ1Rqhm1snSm3eAUcvM3brFnoSsDKac733Qo9KyYWRaMBUC
Etx3v6DwxhxDVAohUnJ3rv5hDSAlWhTuybPMrjVtgdQ7BCtxuiuq9ew+L+AsXgss
QqRToxilUSwvQAjiLd8/oIKZmHF0zU1BpiUUTOcodKdRLTo0CbS46tMKaJx6iIMq
`protect END_PROTECTED
