`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOVemg9SKLNEHzBwuipRIhkHkD1GYJGsgQa9zY9eB7CS
34UnVoSXIYYYzRvuDJSUsrLzF5gQSq9vthijk+ELpaXvqT190AwN5nHwlhJUiuBR
2NT6CsOkSAeDl22BEHPnqhk5aYZmgfpCQUzzQFkYnww=
`protect END_PROTECTED
