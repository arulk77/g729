`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAp8pEW9J+afzQVUO0MeVQtLpQvkIcqNWSRMi2GIo4rG
TEOSbsw6mE2Slq50MXVh1BNeUd90R7YjWsJeAGl9DKqTg83vcgONmI6HnWaljELO
LbU/OWX+Xf6S5Xqu+wZDr+lD5Fy+18Zb0Rf2leMtA0/yfitR/n77wUbm71ykkorC
VqKGC1lvnaEBHWs9wtEbUAC/rDo20kQdGJiMCVyXdVX01GBVNOw1ASSiXhwWQhvE
`protect END_PROTECTED
