`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNVo8VvSZmxJUEUATaaTRY0s0Sy/8aM6MKTHKTd7EX87
2l0SIuCzkef62WsrklkDj39qFB3Hhr3YSXIo5PeKsZ+/cXK5jwA9y6ZuBBOqHtH8
qiJy8GJSLhT5gdycfqwIwBk2NBPU975OL0TaYnbk1z4luEjWFEuI2pgopGMLPRCB
SruYMZ2AaD8WVChMau4zOPjPxfS4T/NoOn5+ycOjJQLFEjWtVPW9Lv0E/FCUwzJH
+TpPYFK71bpr6oSz71UHbGpVCpKjWssm7nJQyH+sRagugxh7ACAwuOJ3gFfbwdzH
+M8S4pIItVD6ED/d6Nbv+VnSdzKFIygos+bn4DoLM+vHQA/95gbPEpsG6vRjCzyU
`protect END_PROTECTED
