`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLbi2l4bgVAwQpfAS+5dNItJljz4pWyTSl2bfBGi/pe2
ErVhxMWPKS/SMvZVzGMqqYm9oqtGuLH7e2hHIvicq6BmbtP00M8PpC9a6DVRgfsk
zsZng7ea7EEmwS6sKBHHTzVvWBfqN9rBr84s8EtkLKxewt/WMW8esJxA7x4xaorE
31mUL8RA8tVUqppbWTuMZg==
`protect END_PROTECTED
