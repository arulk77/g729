`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEgo6rhARQk0RGhhtTKNk2c5fft3i0ptNyx6KYTqfdd4
QmRFHxqwVFu3AxegTc5Hg3kPLomIoUevm+gLLcigXcgqIGPFuACrywk9/xPcNTuG
pZu5NW4UQOWxFZGEWp7PpqMKu37tmIArgp3pS4kpjBHG3qep3THGYMvu+KlvHmxQ
paplzI8x3IrJhnQ4pmwYLA1hOREE9xFpGzqubptkvKH8ghMjZSxkb9eV5XHl2I7A
q6VQHRuSf17QoVxzRr4vE9Kdr0G2wxB5FW42d+ABp3lzUMd1/IPtNi5NEaYSngLt
AJ2SnoPJSYnuczrDBzSPbB/fpebzpBXvEwbybMuNEpgMXQvUszBB6mLOZOOpb2GL
YmQOE6KlOMECe8r+58XEXLkPjISwksc8UQvzMr4t9g1a9EZ6CkV9sTc2JUUgV6gH
zXIk6mVkZhrW8Ue22ZwD1rUSi2rmaq+fnT9jSL+Am4DTzPa2XuT25v2paWueXCBi
eATe8SZY/Cu8w1TJgg9PN2ULrvx/3TxD7PPM71ndduu7aqcA4DJC//MerCpFV9lc
B4eXKQgWp05oQELNSKFFk7m2ULRpyb1GUH6+rEtjUog6TKdu2I96BGoR+0fuzc2q
aP0Qup+Z4tqVn4Z8BAs4xWKBBu1FCkYhzXBYtbLy2WG9C/zT1Lh+Oe2k19cqhXf+
xLIoP7xTqs3ECARqMne0eonTV7YGpkihkzI15LJIqp7OYqD18j44ky4G8kZ7DWW7
QxhBnMoGoq5pRRB34eggjIOq101VRyP4zYsQhVQ6z4NVAhP6ujZSBJrmbCxSf4vO
VcWEUGptSp2n+Rerh1t1/ofHHhZMZVIgEey3V02utMY=
`protect END_PROTECTED
