`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/Q++qJd7+b3q0s+wD75WW7OthAViriNnBo+QaOatTDESVq6PyRp/DQ9FJV+MPV/w
4pKUa+orsza4k5NS/VqplgnbEuNLVfIW5MZALjk5xhlNoo8IbtFp3uk4IBL+/zae
o2RKARNhj40NNQVrYvkvvDDjia8xSIurvzUhqyX4egThYESuwGMEZNdLPT2t2/59
dvjkAsZu2NrNFlt5vDapF8yAlxB1vhaV/KeN9YPQY13Qy21Kc1FeoEfUen3iBLiJ
AK+Bz4ZTfXN9cOrv8RgWYprfhjiFMFjZXBfXVsO3IgpIeeGjGhzSaKNES/3KDR+d
vpKZ3pRkBL4tC5HLmHoZnImKYFrEqhkQNII7LiWhmtlnVtZ3zdnB7ntHNQB3p8El
8wPLAy6Re5MLzK7abslGJ7kUUjF9xBr9xdU3+1RN61/vjLe3CfBRD4OlDI4RZ7Iq
7CsYOkh2hY9U0gEizozoTs964cuBPYClukjt80JBK2jv36kVV7TQF0h72IYvSnON
7mIw6awqeGHLjcpbT15KkuvRJOr0hudG3wBbpOGwabAL4enooJkcummrgdeEFxqN
Uvg6VJsXg5zb/i40qRCa7tVuX9SsQCD8sKqUUHvyN/jCRX36gMy3HRW7nl1TdVAk
vFvnJ6OkPsdEi25YJn43dVIZ/Uvc9Z0jpYyvz1gU0wcnclEnkuKsaLhtL7SWxzjd
4RWuv0Fr1M1LDQeptZHIkOI99sCRmTB/6yFuIjj1XeQVWGVd9oboFRJwd7shmkd6
DdhlUzhRMJr4lmr7/M4ySSoDEPzJif/CpYELlKmHiPwAqgfa/qqhXMx31dVWB2Tc
8173kPctMYhH8EoJDfeK9G5vRuWabbu1rvh03Rr50ThNjVmUmmXKf6GRSzNXhppq
cMjOalJHzEF4T2Hib94pgbbdM8C+OoRALtFcrjFWO5YEiU19+AvRClTHrBKHS+bI
YkFee08J5xXqpgf+qeR7PB/0hOzba/072TswZGI09RyRAwYnxDcvF9XWwzIGW7/a
X6R3hHLFmADD9v3qFakuhDQkV1MTp8FVGS1/DckokGZmqTRuh2xp9dLlNuCZTTcl
llkkSeyeaMJr0oRP+v978XVHAC4m3V/frpHlqP7jsmK+dGlxBRh24nBL99wnS+nq
TfeAgPu0AcqXF3iF3CTZf1Wl5qcT6pMmb4xxspcZSatjQHbEigYZoq/HlgLvmFmi
6Wc66zRrtTAU5AeOK6AScwJnvWTwHDOiaevgbCSJeFu328iHWGAEY/egsors89F1
`protect END_PROTECTED
