`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLfyoV8ukpog2zdoJ664wDRbSAEwyuxL8KLnD9RoCuouW
DO99h91lfZ2hVo8EwP1dmPNKzDEB2O46Z3qXDHFRBubRun0BfeIRiDEe19GqGwg8
tZGs3mMH2hLG6mpyHxeO41FMz7nnpGip1UyTuTuG9KYiTUnzxDyQDHzFtC2Nax42
FRc5n2Ch9l8ZZwddhBcACyHLqenh4DtjfAJYVFC9q+pgMOcHOAbV+xn2ESW73w6O
`protect END_PROTECTED
