`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEbCzHXBvZI/Zfd1Ei3Z9/daC7hmqsi5cmB+sACF/nJ6
j0UqMF4VN+0G5VWHXj4YLNzibOgr5R8kuoke7r4wfS5krTm5YHZQ0I5xcDywrY23
nkP+zu+ymW2zyDzp19r+0ewye8mfBfsil06x/j/xjud7GrAMfwyQk2RxK41DpFNK
TK/iQpwBA0N2wnFIwAu2R/u1FYaKUHhbXxYtwfCWafjIssOrIxKWhWOC6bqE/GrX
wGcP/LAiG3DKv6GeMnlZXycqEHNA0rCm8LBvQHBzZI04A9HEOP1W5UQLdRoEhQht
EdRhGFFlEzr/ZIJyf/moYUP2dC5iGPv+VDQzzjOB5UiOFzMX2zRPHYC5VOnbBs8m
VP749/7hBrsa20XDnTcX0BC0W6VwClun1F9gtHfNKCpb09C2DTyBT1eBavYlDG6W
KI6vnByJ1ASv0CHp6eNKiTDwqGNZvMS8VmeRauOr0xe9tvkxkN3NYiO2RGHH2o3h
n3Gr4qCnafSfKUjD96ofUq6hqQmCUZR+fQJSNy56WR07LG0Sn2KG/HzXGXfPGvgx
+34cW/IYzqI1P+O8CjPOEde/8zm9lmPfVvc2CbH4kReRHn2BvsdjX5FN8FJJ12Ew
J8UW/kz07lupvXA3TAddGS8dwBbobq2vGJ2BROGvcjuXrMSCiSO4QUMO0aqQMB46
`protect END_PROTECTED
