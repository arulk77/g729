`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6X9Z//nw872/ALoCU2+/1MY6l2PCFxJAir+lBB7bSzNec4Jcl4V1ec/xUps1cQUl
gU33DzlopVcXQCL1fuOR1+pAzJqWlksktpLFm8NP1etTldEyKyxHRv9QaN3iGMll
F1VGJAqPwHeokXvvB4Fe2pH7iomobTw5D0sSR3/hh0CHmjluu5QCvbYAS8+djEe7
eZHdJLuOVluUwKbjSg4PDxsR23fgBeUf2d0rj810f3OJYhOXmyVsOvRTXZN6arPj
t92JYROH/wn0ghvUxMjCzf2DUfIhrLVaK5LIByNLbNIDOslBuOgIJ+AWDW+kkDZh
GOCa2R6oXNTYQoofMqqdxllNokoo8dpRByvUKU58iQM=
`protect END_PROTECTED
