`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UPFHi+uh/gFg+9LDlBifND1feAsR2fbFuwxzEb0/yDmx6A5QNW0DMjAxWhp4HUCu
u3tykRvBVKaeslKnngHWWaACR2Wb8sXOMhyOKK2qX/qWpZooPpKK2F3GnVrN/1RJ
uL6I8cZEPnyAtJ08FYD9e4l3XFQgQ0yAI7z4jcIDT9acODSzCyEWRHs9GiKY1ZbD
/WAxODkhpUE15xqB/dAtZkziXI2p2IiuN+svUoL6y/iZkOMUILccMHnpqI5Gd691
duQo46lLogxRHcvG85P/H23PdiYD4GzRY8k3cSsCm0eihrStvVpbLZ5ufT0OlBxL
xrfBCVb/Fx0OowHtchCwGbTWkP/m6P/Ih5sjbgsIKbJtFVsl/+9zWI0p0Q9AOwSJ
vNdjzOvhls30MgoELaFHO9a2W+MujkoPW4Wy1VBRcIc=
`protect END_PROTECTED
