`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN41eJfsXLPBRR2zlrol7TUhJ9HcOmx4YFvxHXhM1/LaQ
/wXXbt0NtyR1hnTHg5PY+1vK+4adpuX6XEWcuzE+qIFuXXvKDXFpis1JMXBRk1Rn
AktxkBFqCJvsZyMeWSkLfi37jgz4Q+40B1sXohto0l7Tf7NED6HlYKAGvFVhJicI
l/+P9R61PtmxRf22ytFLTYL+yyeS87rEkiX1ea76fcmNOgiyzTuyn0a2dN87LuvP
2gVd6VY5Rd87pB/kLgF5njmySK1nQ1lhM6qb5+k0DHnTJ8Fj3bOon/guNpdAx4Mp
IY2QFzkKJnaf3noldpIxeRxIJ2MkpLqgyrbDgYVFaGW4pC45wa203mZ0sgfI4/Ns
GpIhPtUC9P2Kq6YVz77Kv87g6osnBgc9cMnaYoLI00o9E4DKl8LgJFyOziBShaOq
OXqeCRfYh6Zp/kMcnglMyle3rMdpQBnjtEiLzZ+AziZs9x7FHTLsfe9H+8pp/lU5
wnoRgv7TMwqEZoLThoHV/3XRhR1ItKCZYADpmRr+TB68VTs+FEGcYwfUtj1TCvkF
BMDmDHCtxds1qJCzsjZGEH8NoHiUnwsDI3uMlhAlvd8h98Q/wblMmTmxydCUNjph
i7Pk5gxYhVlwMMFIoBpsJvgT28VciGQXbK2LvHdrBlbbSGiV8HXCaGxtPTM334cr
iqVn4iHBLVwVx1qX9DdX8QcQY2F5fAnz0Mnali0RFJKiQAqVphcLyi5ED4Zv8yiw
eA82ttFz0efYD2NwksaLFohx/1BeX4LOHWp4PacfeTOlvIvE9NSuzzy0lI3LS1U2
6lvytr601cP1jTwJuhLvXHeuHqnm2FVnZUwa1cvKrdDynNAPxMyUtJXJ6Cjql3XI
uN4yQT7vrAYOjDGKC8CA/AzaZLtjCORtpLtEoH2/7kWSYXzA8A+qXtUdpNjw9S4Z
kWwftXSWQkMX4PYkBpEuPMODIr950tRysD4wMsILDj33FJqQcLtr4mGNNsq2FwSD
AiuxCrth218sfcPkA+C0pTlPa5+l6qwNc6+un6EnintMJksw/nMZHwYu3rwkd5IL
/7wgt05OddZ+IfRjJO8ojuWzxSNt69XOsLWmzRJAzLWhE2WNj5y+Du+NmUiDZYOe
oaANRuEnzBkMPqo6UAJKEvtlawEqxhJhXF36RGvqhCxNunAENxqK40COEoj0tVVW
RChS2kcNSNpv7L9ApxQJXVBzGc1/975XmeD940Wz9GzPPmWTFFMTKydpZoLSds8t
2UGPanYDhmXjNrRKP4mBVBLtB0CouQcct+u8uxJtCBbUs3ZHc5dCcGBDPVVDuO0f
hUxDL4/Pt5FjvyvkMfeYKmYOzHGexvSqVyjpmUKecP0BD/xiHBOeS/q3AARqQyc7
YKc1aKyGJzi5DsAPHje7nMJ/AS9qKBaA9vbyk1s5Bx7F1UsXsO8QtI41T/I5E5TS
FcN9wk27bXFTiigphuTCp1fg8SqG6oDyCwnGOlY8woktkYS1Tv1IZrVAs/EDDMyW
14iBI83Mq/DldNmKargi6tA0VDE2OkfsM3uWqL/z/BGXf+qEMMIJGbNzHf5y5q1x
I6chAfF2qQ2YTlnQ3wuKahCsuUFUA6tmfkxAtWrA1T7xPDmDIAc0CIOz4W0LA2Xy
xgaFdIeW5IdAeUQjb0uQNhAP/wvDLbyHXDTCgQAwnvBquR31bqOwO9CiUC/tzrBC
kwLhi/xMIlUBRNFn4rSF5o0UrKoB8dLLka9OMjwKJN1rfzcRWRNUj/4IpfqErz+Y
XqnBmPA6OSo/4gSkliqP+YXFKLOZCq5CyS3wPdDiFd8x2BqMVQxJQFydStAeBr3b
5+6QK1MPxxy6WTvEYWxC/Cgc/2vQ6VDAzM6PxtpL6ln57yPQcyLBhAygQsZpMH2G
zK+iWHGIFcqlNief9vDr1vk75NSiPN+imPcLa1lqXED3o/8kUHg6Xjx4M5mf53Mw
C5D8/S1LXs/OOB6CwSRIvPwyOLAJ63oWPIL9bZxXGezagx8BO17Lt7p0YKN0QgcF
iJaeAy9bKY5MHcEQSuqRHisihHRnZO8PF3wwxMT3Mqt1VyyQt3Yea+fSV7s1cv0k
I3pRSw09yqgyftkzo0rRlM8IfX3fQPXdJonxFiTBUaoTAK04hPUxUuVsZDELb9UZ
AY/RtZ6OWlDarxa6Cfi1WG+w4PkDDxzYeGuJbO/UVVOwShNa3H9UfniTtz2XZp64
lXIxHHKR1XFbomjGnOq9CIPz0uRPwAzhaOe/Yp3uY6qkP1Yp4Y0FUW6jxsDg4rkO
i7VyhGf1SsepUBJfrvklW2XFC0whDa/wqzw9EUopcBiNQica0WtDH2seskEMdIfL
Lu9Dis1wUTOSoPxVvlXGXAGHRdw/dw0bythm4vsuOB9UVfb2+8vpmXSDLuYFW2ux
qs5HLkw5mUSvBwg1lw6H1l8XLDV/SxXpN6+AS4/uO/VNJHWruDmIF0KS7EpWEv+t
0OQjficmR7IGu832XSemnbTVt6TJoOyjsIIWJbKRgIZSuIUNYNIccsWgld9YS6HQ
kRYFji6OqgZmrF6gvxwPZ6sfRW51omNjhJXeIbP5hWqhmQOCvpDKeaHfJTKFO0uF
4yCGpK1rGSCYYgGz+Mbz83SAFnBORp3PeL4yU4HPiyHbnKK1Fd21uKmlafl7zYiT
/4gSPCpdopUcxyA8NrpJggwuZmsdiLpyn5J/WfROKXi4Y39rxgXyXEdvDB8DhLUc
h7jWoAZmHDL9WBeNCPFsWf+hWFICbZG6me8y1X+ZOLq6BEs2sHqLUkNAc5lvolji
9FoUfQTPAjmWpy4DcbOac4846Yw0N8jGMAOnibLpfCmlBzkbJW54QekY7C3vrQuf
DhVmKGj5ofe58vwO6NCkdO8kz9Vi92sR3LHPoBma65XuY6xaGu2kCjUeKSco44ud
P7dLrSd64mkQEejpMVxnSrH4SQtn4PO3hyd3b3UWaepQ+lpo6HnvVcqCdEBmCSql
QYxcnnGqIlPaF+y9O1FO8ftHMkWcyIKDz1S/JngaW4dLCBxmdcBM4XW5qT4rbW96
1T1SHjMA+Vu4i2NbFU/Z2wW06C6AxtGgzXzS1WC3d2rDwZW3pxXLzokGCiCUDGK6
TXCv74ZcLnqtif9fToy/vxP/ed8JL8kYuJtQoWjyiM7G6mAfQYKDLZLMb6+8VUsr
/0vinx7MhmJOFtw5uagb6limIbfwgfuNP1rNWr9i56Ikv1yPxXZVBCqxFzFKUXRW
xYd/2ERGxUQXiBzsdkxtT91kGeCRnGLIIWgE0zUk/3R2yUfFPjndMF0VJh5lzrR+
5gpEPsYl/IbhFB7t1kDw3il5Hbuw8Ol27+iWCLAjbcXfCVpGfPdWOonpcN0Fb524
WJD1XXyI5WXbx37Lq7p8tJmoS21GMYpG4+LLjWl0WbqmAUR3qECCw9XIZeR1Gz3j
pTpZ6AEwIaKW5sdMQmMctwdpOH3PuaIcYm+TNMLNEpTTSwpO072CWK+BxUbDxF2M
sSggPRGZ8tcnUA9awj5L0pGLDTShMl3p0Nr4x3dqhmcJePuieVkKvDCPFAUAim4a
P4swtL7jjD7Wnufo4i4aUkW/qTq+fxXLoVjtFJxKpCaQLgQfVOSKiHmgSDp9gaKE
m1xPDR1teMnmbQbJqJhx4T/4v1DkaCRLqcrzn+1x6qCSRRu9heLEOQTG7zlkL8I1
qO3vP9x11LA4SsnGALiSlWGGGF0nZXy8BfWHFUKnTVnXjRCQRDA7RoayyX05nCME
0fU0HWYSwopdRS2PCktyfUi47YbC2/1wSszU8Ujj77V57dNQDtvO1NdvtZEaY0B2
V4ooYbBAbtu0mFPHVLJ3k9ThKbJleXhXIIgP44Z8IpOobFH9RZ/cJiQ+B5doY4r1
9h6Eke3wvHWWeVWeIFez1JONAcZP1a97a8yVv3T7OocVvJtW8AOdFCb5e3gwCHAy
xuV6dHZd41Jo8weS7cFpq2P+Wd6dWml5v70XVckvCC9ojK1thlhTMyu4bMXcNSY3
CmRBcaSRV+3whOsq2fKl4TE1mcx8NsTrHB4hwpOq411XOJWxPTsQ4M/VOfgTzIdO
XMZQ3Erhqoj/2SUFpgDBYk/g1mF+mpxyLXpURzObe//HnoOC6MoOrzqXXO/4+gFa
M0TDNvweSxg18niJejCGsZMpJ3QtRwni8w5a78odBA1AyHWkuxxoHu/0J2w6w9ma
hXRG3nbfL7led9kO1TQP/OrmEb3YmNmNoYN40HyajO7Ve4XlQ72XiCLpX5yTMoGe
VYevrRlsCBvEMbHOvoKDbhuQaoCofJHKMpY60rLdNxD6dfLWxrBOapumjO/shAG6
jwKluGRQdfN9IEZUNmn4YUnSL3yEl7mpUPD4YLJEYMLauJW7CJBIXVoY3GxLoVNu
nBS7IXHjYMv5wiecPeRPBZVHsQR6eZ0dSYRgC6KX6ofjIEahNmfTEfX6mPJUfO0c
wQ/nohPJPqrUU0PonMsEqMzkYkytAKmiZdMK7XZGxXVE9x2Il7eDj394XENSfJqZ
9bR9KyhZ89hhEfMtenkpSNBrKYYBLVzSKJLxOcFlnltgxTjsD5ZcQ2MRumWAwDf5
kGgn2+TH7et/l+CG3PjfCGddTzfoxTgWn9HpyxQopt4SvA/a50JqvlAKBO12hDvR
aA5KV8AW5C/4seLW1DMztColTxeQuct46bvZeFlkFEeqMGtHCejvm2GYcHmqt4SB
tG0ykmN48MzkIMeRnU1mJBE016MA0OBycrlkiD7FE7CdLe9XtcfP1iXVBF7s/E49
W0HyRUC0UQhUWL0ayRTk0yF4oZnvy0skQoQYnpFT4RkDkGOhrrXyQaVx1rXLnXAD
mti6Kfci+OyAzWn+5W2r5R/Ta8iAdv9e2dc2rldK9VIxyFoCyAiLuof/Joy8aZXS
5pPYvDQ9GJ+4OdoTdvTiXM06raCUm+G6TPnyf3kUP+N42Fno85RQm2QZTbnK/Eth
8uKlfoZ2LXcOkZ+BWsViY2oJtf96V3YxDWNfw52hY016XlLri0/rfsQY4Q+gnEMN
AQnWtDi26qH1rhFyW9a9szO7wuip/ps15BjMGaXpkL+Ibj6+LTjh0gVxBMICG/zC
UOkHgGBvQsSQS4tPnibSJ6WhbdYuEwQXYu7NtEX42EHV/nUiI7qSg2JObveBsFrC
TJha6o/3E/bfzKEGyC6Bc+VelkOCFE5ifHDzxAB78HHiXiHe6VbxAO9cdUMbev4Z
FHoEC1sgd7NdChEEW42CYRI6FftWThtgUPgYdCouWEB/TuAkf7lEU9vRhI+QEPdA
q2SozfcWGLBgfDaSaLXPuZWHvWwrEz+JWVJApfCkW9JNcDxRjcA8zQYWkdQGoWHO
7xZ/12YPNa+IQNgLQ28Z3c9YJ5Kk+wuhMA833jQiVDTzkN8UYtR0TytvWM5PDPRe
iupHlkcZfT4UDuE7vAMCUkvbP79zMKiYtmXYYuWIK+SQmN0z1SH4+exrn6opH7WJ
F+xF0szDbNlbJbait8oBlp2NfOXEHgAHQ4ItSWhMuTvQoGAQoO+McKz0BLVd76K1
AGkdLEenCY1yrNhGZUBIjTektYU0OK0c5RcPFKnPYC9FhuBDJ2dXnRNwnZK9WCQx
QtSwpTyu7a6R+a9otR6IISB+viRcN7x5arOX+/W73yESBk+Uw+Vop2Tb+721VBcE
lIm4XqY1MUGuPIq58ZmkVHjctQGA8NNQIAktxKH/nxC3J29GKTOGBgg6eHBlPnR2
kzSfkyZPM55McMT+k/Cyq5488ef4SF6wWeRZH4T2HKmBS7EAJh0wWyt73ZJbh7l9
arlQDMFSyzc0nH0tDPbhshco3NUWRZqauNNoVotexCYYshv+BDouuQ68Mk1J8cXH
8OyNzqJqkWUO3wsROxcLp0TLfj54o/D4nkRKKlzw52nYHBWVQqLSE25x+kjajswn
8149RfO04Qk24t91FGJych/rz+SjTiIyMC6IzeDPuV+xVrKejeAUD3WSpQGVIgN3
YpqLq733QXtAmnUJ0lutKIyFzpMkmsXi5jTxhKC9r987bFjCSsQLei+2dq+q090v
0DphHAPP8U653uL1p5zybR4YNe1rjhT3sFSrjz5vrpdkDTYeqa+m0cRrnRXjo1L7
6xw5dBsu8g5oKCP6JcL4GTytsPsm04c1vfNwtf4auVfj6F0N75Q8NSUPaxgPUJ/z
ptsHx/0n0qAZcR9qWBZICmTdaJXaq3hk8QU078/YVSCEXceJ/VfMpakP8QEIM+ys
wK0OG+YLghCqfJgSyS4C5yjACYie28VAo4t0p5MC3rYQY4PQglR6Iunp+tbNOQ9U
eR2td/kL9LJti9jn5sEkgoPnN2v9WV/OKKzhtnrCjEbSJqdFKkWHDIBoI/Lu+qHp
9Bj7bplDjNkSdcbGVKA92OGQ7la/1+sIzuwpgupVGFrkntBnKMVTSzzF2j7kmnB3
TC+GNTotTiX7G1fqD1UzxX8ClZe9Am/XM8mEWYRLELwTUtG/X4eC3kSjkehi8f9+
pZqmOwHNK++BSCKOJQ5YKdXsPSIz0SnXNcdfjgabe+iqVqZRrgqDuoAswWqYdget
e9AXwzsHCS0U1JToqWBYtP6K2fXA171qBXwQWDXRxejz3Y6bCAw5aDxzL/i62+0w
PhztvS3HTsTelUm6KNh4p7A0ZCbIhaue1Ua1xP0TA1bgd88WJm45eB15QI8uSrcs
fKZ8+i7+lAFIds5gkmo4dS6ka72VSMMiQFp9sZY/T1IORAAL7GALrWN58yoIUlBC
`protect END_PROTECTED
