`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGrJDfWfMeu199ZFZgg3sYSLpiqtpBoHdrM3JovQK8hK
9F/Z/n8nOeOLJ1gE9aao5jj66MY44P6FNreFEmlrPdqg0ayMrBDMfyidAw6TrvF/
6phHWUT2ngJjmwRMOWfzyhU1dga78GLWsZ3moHjjd4ziW6UPvwLERvcyJXhKZ8Wq
x0IRxTOeX0LTf/zxf7XNudv7ajZ5fgOBpg8DBHfVI+P9j0sWGhHQmspOhvmXbz0Z
`protect END_PROTECTED
