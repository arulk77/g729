`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ePPHfYRSEICaOLoLN7FVu62OZMO0hB24U/s4vth0pkU61y0/C174MjhxwdjePott
imo5gGx0UDbDqc/w9QHjw3Qs2yCgWmfbNLoHc5GkAZK3tcqEHXQarqrvQqFFJThq
EQaVHSgf8Ci1+hCBAeTtZvF+/ZZGIVkzSmkP1n4KW9b/Nh3mUz0z8A2YgLb9fMUS
semxG0J38wKQYPtCHaIdAkQiyBwqUWacWNYTahwlPikq8KNfCn8plQWHQDR3UEpp
`protect END_PROTECTED
