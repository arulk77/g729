`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMGObKO3b9W800TS3YcQ7iqFJJ0hyYg3FnupxnpG2hEE
2f1IcL2olAYNkAfsdJbmTEuq5k5+DhAdGhfWhX3f/Ms7Z7vBlVJ6cZYKCkpb5pjT
gyDcEurHbsgNQ386CM/GcQFejiT8fVWbIWfE6vnplb7IQVCNtIvo2yeMu/CFPJ1N
bSJzoeJ9AW6GqUddg0s+uSLzIbyLTZjTGH70luXG6CNuqVR0cMAaerxYHamlugJa
HWioRd3dxIimYKXbVvkiVE+R5eLRJ4aqD7qPPhKZ0wkco75Hcw91MFRjOVvzMPwZ
VgtAIKl636b3TYSnVECoNpzPNww2gMlo99IKx1IUoVZNzylAeLzEmol7DAvfiZAs
2eKjZhovN3y+fKf3bve45ZMK+BIOUEvngL4ix06xWNjAeK5DCaD80bVcdyDZ4Oyf
`protect END_PROTECTED
