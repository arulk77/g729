`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveChoSs+CrWyo/hwLtHfqx6AFfLT6nYLmnjYNSol5K9nT
KAH0U+Rp8sSElGjgRFWjYWt8CtitNR/4qq4XQnKKddjYjiwb4Ek00taACSHo0yDI
J9YL2FduwxJSmnMvMIPVKQYZE8quGeGqkGWtOMIxN3sv/NtOR6mTOLNuuMNn4jRz
NlKa6Ic7RgKwek59u8ydUA+xBEr5OFNePsuhePGJjdez0cyoAEdUjwEPoVNeldM5
ONgtWSGI90lWQok2fPYGrDPS8wp00iB+OSYq+qg/KdvKTvpTeDtHv/k7eDgm93s+
owaSq0jKIKORlZF0n0+Fr5EuZBJNtknFvUT2AyUwuY+auFUMjAMCAvs6QAydy6MZ
PBKLei3KVGnNADfUM9cSTPyCob06VnvmXFSkXDDnxbJlBlCv0jDLGQ1wHdzpSNQL
z/gSY0rzFyacB1bPiIxPe/15uSjhQXd1Tb4Fu01j4GW/TfjGgsdSNT6BfBY6JSNQ
Gn6WG79Dsc0cAl8+RtO+8A==
`protect END_PROTECTED
