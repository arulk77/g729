`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40X8l6e7P6sUhFIES0dbe3e5BBlPEgceIo+OT2Ws610x
Hjert7UQ4D5EvIrNA46qpIJ2jgoztOQzCTmvcrGUiXyg0W+SVVSc9O3crpoA6+Zw
RkpKp7H/LCtwOylq8MFngy2UnVfybyTeaWrhdpp6u64XzjxRkQ/uIESduXhbqZx/
bYIK8X/IkdiRQuMq0bGvgJWH8iFMt4Rf/Ve4mmAld4lO22tk4nAYoAPg0QExILRk
cQ0tUFhWw8PsqYzA1RjzD7DspHxLdxh6wEWkyJG149I=
`protect END_PROTECTED
