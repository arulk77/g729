`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIV3M/0PJxNx6mGQj/ZgLAAFlzXhoi0D+JnN3g1OFj1w
rssko6BRo8PrpW9mkmVKsZ4MnT62YVWaa2zrrFdEZkHuL+Vj6RHvWFJzUiRpdCiW
RSknFUbCRGIvcGGPwr9zvbvZBFyKlqpFq94eviD6z2fscD1v/kd5KqZK6sHd0iBu
fmQwyKr0axWhbXPAKSXNGA==
`protect END_PROTECTED
