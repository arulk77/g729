`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
G6kA8ivcKGk04MMHgK/a313Bw1+sho97nkBwqvAD9jQ5RexvHsaZSGkQsVuu+kBW
0N6ewxO5cW9mnkO+mQQ3n93AnCnVtCgJJhuMAnfdAO4ghs8d8OiDuVWFQtBcEPPy
Be0Wb9tXl9sqK3xoN7jea1Pyb8uBBEPuJV59z1AXjI5hjaHQ7WMf+QSRqDLWRwvR
9mvvls92IMVnZbJANs5Yd9zNtWL0V7mcR7GGr1ubXfahC9lUHqHoJGmgYRLaS1O+
Ud5BOHECnlRSotcBmJegy33gZklPmNVQ+TMEYA2DXz4=
`protect END_PROTECTED
