`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
A+ZrOxrfe/NWFU4TitY2st5rBLZa2KJCCuKSrX7Bqu3EHcyUf+S5W9BVG4uuLx3E
4XifJBxnb2zbiBKANGUxhT8DQu9Hgi1Os1oVRnWcjIaEhkTbyGI3c5obOilVKOme
uSpyzk1NZSWvGsXdQA3z+elnNRfjAQrpL8aDjvOX2rTbXaJwf6mHDbBgSYpR8J6B
vaf9DmupVQ+ZutLLLEwGszB/iBdOEJWhAdJ03/LvuL8SBI+bxJwXpk8G/u/PT71A
DK7KiREwoYF67HYYkgxiXnuxl6xEXAQssxTdVyjdCCA=
`protect END_PROTECTED
