`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHzLMHobSAmtMpwEeW5b8FT6Rwu/NTRy3awz0ZiFE2GU
Hwi5gQ7NYtXsYdbg+kBcPv5hu+wlcJnSnxKd2al6uBpyyXE671GsmCanbRpIBDBw
oivqGCoU1YeVeZY3T3KkxP0GyzcBxgXcX20uv4iqVNImQszjZTTXZz41zaqcW1dM
+puWkPJMZLgfo2X3ieEyVNpd6WpQ5/6r7dKq4U6X518A6e3qKHLz+XX4l897OB5j
XmdSgs4ilSVZbH/cqQDy8vTyi62HOBqF11FokgvwAA1UsknVlGFVCqwnB9pwJEeH
jimrNOXUlM6hBe0nqEJ53VBCo0uTUEzMNoJbkVEHvKLZ3RgW5fO6qIg/FGxpp2Za
hXXoV7MbrFVgCOEv48qwR+GxHJ5X+HOU2bHV78M+5oeemuBdClRPslWVSL1nTCMp
Fa4InwGCB1cEy5zg4Pt6Kk5HZlSSn3cZV0wmLwn1nnAvju4Bgs1qzmtbIaMJ++d1
Onxs1lGUaHbtpq+yn2hSD8tTuSWQcJ1Jz59SGpwvx+UlI2tIbiEvxcKvwNFa1a4+
vAk2rNRUO/nUB+1hM244mA==
`protect END_PROTECTED
