`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu447BIFft6YnWEpVCyUh9VUvEKcTAtRdVUFnbpIJ1KxsW
NzodxoeqbyMa7wHz79cJLPnxftKlzkcwqCCj+1NWRG+OfOv9RHvfzoxtz4VSfeHD
C5yARn8zhVisAJ1gMcBKLM0XG7bub8xxb+SumqS1R65p5X8sM8FcDKIxAL3hlEGi
gN2CN8OvTcbD8N+cxdhaotqcug8n2+VfXzKe3lkSmlPMeX0OdXC/2HVxuUC7wxS5
uq/olb0zRvEAvwRE59zm+O+t5RaI24TXAei9DVrDZa0=
`protect END_PROTECTED
