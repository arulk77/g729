`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
R2KBd7yoOiQJtLLJH4faNytNeBQ+ocyi3kkHxgg4O4+Cz9AqVO6e5bLDXchZiYdy
29tp3GBXoMNaO9HH0vSgjHdQ5LKLoRhIx6DI9Pk3K2Ey5n+hlz6GqRmV5v8djbwi
tKBmPZQeLnYbEf+HoED6wQiztzlnYrpPuGAquank+Mkvp3cZAU9Cdio72mAJEEx3
1of/MTuYZedXwnO2v24rjZhaCbozuZSpQSNNmuBKeirDats6+ZE28S7qyAEPmYiu
`protect END_PROTECTED
