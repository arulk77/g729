`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47FixqmlJ/jDKztQ+cqvxuHupWCkks/+oSUIlmVyV31q
jeyJB3cKjTl74xfpceOCfim7qVIZ+9YG07Y4NcA0ZQYB2v4HBM0TSr2FVVq2iOLi
4SqfO8SjnYg85s1A/NVa/akUunqd+EURn4yZSl4+Hxcf26NEh6dHFQCCClfdm6+4
nkJ0454iIAzsAf/AMBgGi1GVg+YrbWc5x2FAKCPJqSXH6ICTrBuDChEb4mxSYwli
pzy+qsMe2jNborknLFeT22DoW5TsM99NG6EIubVeby4m6M14wCerxqJZtpIruDi2
5unWep8XN41dD+JaNPUY/wSvuEBWAHo75u42vXwUsSB7+31CtuS5LdHNumSUsFIV
lzmK1VMFm2tyoMzT9Bc2mQ==
`protect END_PROTECTED
