`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxTbUEntawsTi0c/147TdgsEAlvWonqC8jAWHesLP/4H
tiNOwVSSycR0ZBa0DYL47jdIjiIH8vCZ92GXKQVxk5k0yxhwJm1Mfv4Iq5rVekqj
xGhv3Bu3N+CxcAQMmbfGKrwbR6xw2d/4QB9HJSniWVPicXF7XwXbxn7WCCiLmzZH
AsyYcGk4JrY8OcAlkEc863zTFZYY/xPapUtwhMCc2/iQpuxnVueJ69/2n/Ie9SAg
dLOedOgSO/GkQIbpIh76W3oR/58wlfBvuwwSDyZKh8Rb6CyDZJkR1N3CsNZzUSry
7/FzDRcnbjZgWau8KJ1WuDyrGWAvsw3fKGdBHap/5EfFnoagPKGVE94QMFm1g68A
Wninzpsqtm1iiGhvcIij/EPMru5VadbNO3FtpD0zdv43I6oIaDZDjfBN1lkNVoGM
EFrxkG8hIW+NmRAWCOgFaOSWQdPqmRdbsN17pxfa0wZHuSfWt6QUmGIpeOHOfOLn
UgBlKg3l73HzYpfQHOfVKLpG9OX0t3B38DNOuhAbl4XLXv2BYmDbdQU06KhG2KGD
YaCO5SnvQE+eZIo1qyqddeXOta3L+zrURsmoTxDXIGUS7qEMxI4vSJqd/Wigpqxp
nMioGkNaVKC2Rp9xEN9fhw==
`protect END_PROTECTED
