`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GlKNyXNm+yZpZedmpVG97gcSf5YLf3oH8SP3GUR+0MXj/aP3ZMRkrxzC+j2N6ch/
TAOjftrkNgDouSfHiuT8/+vPngb1pnz0YobyF1tTCesJrKSmEMPTws35DI4gftF0
2PvELKjFPKM+yd/WUBIwFw6pmymrNh3buJZp2zls2GJ42wqmUDzM6TsmMuTR0ryP
vFrBGdPxTHc1cEWA3b4+yYUI3Jq3qYR1cg3fzfpcHyL/EWf+/JBj/NWexpJFrYko
U2yZNM98+Uu99zSUuoOwH+z4nhd5lQQww+Cw0/ESdiDrIrEoHNjosN9WzCV9dwpW
pHnFwK3RCx+B+uAra3LSArpEZRA/oTeCH4osLmmxltT+G8wF9Jg5viL7sllwnZlD
GymyWjLOYf+dppvEKujEyGFThFThd33YVgPRHUb3z/kLT3P//Yhgul8bbhWZMzwx
+ih4MGp+Zsq2Kn4QrwSyCPsXiE3SClcn7rrR36q4ML5tUZGx0zIalbFSJe4ajDx/
GWgacq3fm8AtSyTYjAmFnOMYqNA9DemPSAnTGyyqSNHQXiWzE5mwGeYF1TklAaJG
YwVvDkBAI6FWFNhQmNrdHA==
`protect END_PROTECTED
