`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNzl6Hrt0+VT9Qwd5waC80mgnpZd0a7kpiMjVlPCYr7Id
/JKgRWuAXoCdAv0XYvbvZJ5KOMa4mFi7c/Po4MPBQ8YcCOvJPHOZQ4zjuce7j1/a
VPUf3HEq1OGbfFl0KPt96TchiDEb4q/m9D1ZaSDPSE7RdHBBg7mA3dWTCX14EQRx
rPcr1QM1NZ9UxvS7sP676wwkZD0GvzS6ySqF31VFp3ZPqZCO6S/DZ0BfV7W6SNsI
B6o609GOhO40uhXGbM6XzI9UbcTiaXHTrLxgLScfanCLKsyQPOe5NCadlvlBHr1/
ugmO/u+DSdow31O/jjv/DRUqbFYFYJmUMt1jcsp61x7ohdRg0EKvenIwfvLVJoWJ
IQgVl21fiPSNPl9etp6n9lspMOzsfz+aK6Gk0UbeywVdR03zs99Ogkqb3FivRUkq
T+uivjdEc4PzgzOX4tz4yNIlWJxqhkfz921mH3qoBgsoaT2a5cVFJWM/C2O8qt15
2+RA5EmrQU4RzrUm6t2LoiUDqC1RaWWTyX+DS7KbkEe0MjIf7vxTbq1/PtZpbmUg
5bsH2UzCbPgSQA8iXaxTlKb8ezObd0id9x6+Ri4EDkwCpWY0Kyon8XAqjxJ7sUZv
j4dIVRGrCr2iyMGIiZvB18iUGReNTXAhyyWjhHIeGiZVnSTIckfEXFWF0o5Uh2mD
/GQmRNF5QSv4bcM+1Z90H7rscuu95G0/hVwrxENQRASIpfwkq60qi1MElWDnvEct
RydUlW0d4a8HRqVaJN+pV6HBN7jPANCeNsdRpsbj39kQfGiFnCBOjpYrlXAbrD8u
W9vAOcLw4fiB8Uv+oKaRCDUxtWiGs9/N/ZGE6bnVW0mOJSvazTOLBVoVUABTDMWn
0G8sAJqVgK/jgMnycchu2DrBNmNDu2CIu+gx+pbWLTAvcnhdHONWO4/Vjef3cHBO
hX4WZRZjGeF91x5VCWCjcNLl5hzoyV6BZ8LDIhF5QmY=
`protect END_PROTECTED
