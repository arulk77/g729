`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH6+bgj/icWRUv1u+SY6RCUlsH6XAqwkfg0gTGOppWSr
jbWk3/M7PCkAehJByplNVsQe2naHkE8bdNIfTI+LTDHAJClBPIa6E7hVPIROi6n7
Pus3Wj+4DFPImN+GAO4iofy5nFMJtAMPjcoJlYEFYk3ZB+X2ptkq9O7cXjfkauD/
SQg31F2NwEx85YRBM0wzPIqMk2C0f2Gc+6kRBPm3F8ATdwtftVHH3Inelv+stZCX
gl3OaQsxYlvPwS9g38IqS27q4QJshEvLOwk1wD8OXQMXeHLmIarIlRyCu6X3PCRY
Y93RVfOCWQ4K+k7yGjJCizr/UBkpnimxaaV34XGqNWZ9Kwn9qaNJvoSaeyfW+8WZ
c+T1ruYauJZ675iMg5MoAw==
`protect END_PROTECTED
