`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFE57pNmf5Nykwwo/+eN0Q//SeT6Y+W5Q8WP9IDgpDAF
qoWLuKiuOx76ZBG0TgPnilKpwuaIGpbzcvxl0nyhdRsxeIugttcrt1Z0u4vgcK4Q
OgZL7LgO8pQY2blYNimRGvgED/+zlN2LQMG71dkiK3uaXUPGhbxLRLy6Pstnhi3n
M+Y+ciIxy6ue0Uw6LYe0aw1SkQ+AqADwmGqYXVw4sxdXp1PgmblnCOMXufaVe2je
`protect END_PROTECTED
