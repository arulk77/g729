`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
I3dYFhfxSoyEGJ51LMWZlSuNJwpbmHABoLx9vUXu/Xczy6CmYP6D6SI/3yKkfCGC
0p4PXxauA/zNccI/sF5ParcOJImntFnjE6d+4on+HZNlOWKq1bOjK+ZvlhGon2DH
jOiddyJNIFhhE5feIvPD+uewMNnQaJqT/QnRBg4+WjbwBSN1Y2Sdccrjh5Zvdppk
hw+Ssx+04tviBfEqx7ldeT497zBqQMurza40r6r9eUgbROu0nQJ42NlJxYKfaZC/
phGOUYRm1Z4lo/zIbsVQYg2oI5SGusu5TC+kALM3jrrIACSrB++ALFw9vkG8V1m4
yPmXfPng+dYi/FiyAR4FsFz6lC1RPPiXlpRaO+du1Bk=
`protect END_PROTECTED
