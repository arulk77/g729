`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDIWh8nLcrYH/MkW2lFdVWJsB0yOwf5bOrc2Eqjuk/4P
VPrXfylpZKCuKUHg7axG0c3kmCYvc20fS1+KrCgLOoPdY2YmxyV7nr4wRe5GxUlE
O/BB7ujarqb7h80WqJHIOzYre4Paorj7aJs71vS9DnOUDL67cfqb/t5pIVmINfRL
p00T7nZbk6OJgQCimbXsb+itnhmJNvAdMolIKEBweRc6nQ16Sx/0TAOUwUQquy1k
DGyMqWKRSc39Rj+f0Qf5imX0Qt1KRDtqm/oW9v2/zJNBRIP3ctuKUAR54c0baYPb
j1sTp+QfzvBQVYUB+CETy2dDTLwNHtpVwYQDczaC7NNGJ2FwCRxCKhtCjFx5BThH
l8Oduktn11aOThyaHRrmRrET/VTTXilaGquOgWuQOb6UcGwe6hvP0smmKay+I1XS
S8wwqCcWemoFmxWZf7vpdJxnNv5GCJbCZxFOgC3kOIxDZ0W+fimoDQEGhHD5VBzb
`protect END_PROTECTED
