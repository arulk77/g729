`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xNLrtmhMWddBnA3sGKUyvbrhZZHApwy5kV2sT+cgofL
H90dSpQPXWH1Y5i/QOcV+rgK3Sf7r9mj94M+Eit044l/Hfmsw8etn2aH6eN+Ak81
LMQwq035phiTeqj5PelTi/9mBFcHnmCRZC2FiPS3YFmqAvO0NdFOWgMhcTwlwD81
wPMxoDTiIEJ1qG1l/OwacLGqb1VOsIOyyfBWG00B9PN+69Yb52hpd03C+7IeAura
7e9ZwoMJtva1ncHOqjaoCVb8lDWXgwknrIWRKQEUtPxSWAWgnL5vrEQV2lOKQRb4
PQGesrTkXRAG8sVWz2O6ow==
`protect END_PROTECTED
