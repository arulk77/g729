`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBxYl5W+99Q8kMzLEPIAFVWX+sgUHa6eQWRXO2Xf5+fl
zqOZUpaKH0onjpDjaWoBr3+m18pZZHy0k1/LbXZRn+bg/ke6hVlX3nAbz++XWtUi
8cr2SxYvxCIaJgOYNtToU20cv4lKl8UclsmM6XsosFEeNZhTX3d0A9yBQm4S/VkB
vGjzNk1qpetSP5S3NxTrI9O7BZaSoP5PcLqiJbo6t/yyt/hobScNgLqnXgzlLlip
nIuyoIEAgJ9iyAiG4oYNn47Xvh0ybWvd4f9g4k/4NNoWBgIFyikwisfkMla5YoSC
VDOMq4DoGM36DUZqasP974m+YER4E7ivw/jWyipOijixZ895q0p9Cuw/U1DzmkLS
I9TYV15oRmA0Emr+oHX8JA==
`protect END_PROTECTED
