`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SebokVCrhvG0//WmqIIz93ZM+lZAhr4jL/TAHO6HHieG
EDbo9OzoGdKDf5PiPzZFjaYNzOA/aFlF0jE7vg2F5f/MVnYV9vlC+sWTbpvttehL
PCzYVihC2L/XYxiKsIfG9uqWMDlRpgoQId6jiwFZ1cV+9u96Li0xNF90OA1flYh7
fjId1wHvS118rwaVmHXnlxcUkDFcFi8QO40ubpvsuoj1/VJrwGR1nEpZJOHK0390
vkSCA3ilWbovbGcyAD+e2nNRyc6HSNta5tTl17D4T2fi7JlkiLFrktVPXqOikVtN
CaNEpSUNfciNPdCZH2d/ND4y4ErnphX/OP3IWjIA4f5LtRBImjibMb7MRyFEaOGw
N4jlZJh83IfLg3/As+uXciZnL3xW5tMjaNG7iecV7Cu+FkCTRlyqQMMtQHBKVHWa
IBNRcDjpNp8PKvvvuWro+B1StGAUott2PxODGv5evi6FRTYs1/DSNNEUF5v3lLa4
RPLPd0Y9+myntl6IHn2M3IQXkJZSSSgPdgWpiBsQBDTL+l9a/EZRCrFEcYOpXxhR
Hv/lXNDV3/i9q0pW2n2QpOTILN4QXZbWYEcAMWyBRft/jwFux1nKiUr7J1sef38i
874qAkqUYVzjH+TRcLhA9Ijm43uJ03kzL/VyPOXLWal1iKz50S9tKzDPinm+vbVa
hlUsmz+njdpm35b8RVz3clMBkaniD1Bz8mWGxFfURcmFhr62N3H/8bX0Q4TSDNkk
jfpryFlxjidGmylCAO4PquOe+EKhVSDkmn1HxaxDJOiDoiTT+79o58IP68UznS1j
d33tTC5DK4doxcRZqiXopTR8MFWmVNll0K66+RCKIwmx1rhRYdbXXGgBJM1MKaHq
KnACjmKE3SxBhdFla6GRDDMjn7Ap9MCPGHBTjR7KJCanFL8qrf/WdXJyBbntP+g8
0h+ey2C0vPmnlYbKn/ePkx3SvIWWdJpN22AJW2Evhd1NooAdUfRRQaWegcsNsllZ
aMHc7YGIy31Bm+TnfUMpfx/1TWPxACzVnsfA7YVSQ94mkXsA7I3RsDWtWXhoJi5e
WJ8jT+SUHVWTq/uuBj2KsDO44fYKAizNHP4BL0IE7IB+qn8QCV5ztIH+MrT8LNcH
g2bIXgUfu9tUjGLJNuWrtr8IVjXvVJygRa5HR5VDt3eQPSNc/l/w4iu0xE3DQzTP
v3bZIuYVoctQD0/AU1+CzSRPe1KRa/vCBi/c1TdFXsH1FOPTeNB2jopFNwpKAaTR
2A4Iy0XfcJNMGeA4J748KFk2yaKEL2Y36FpgNOkwRycQo/2C171OLGbQOMkCdSeH
VlYgGOXpU9DW1ZJ9GZzHrCQh0LdKfYShDqoCdwrtN34E5/Xrg6M82tMEtLGAbrmy
f2CdEdnwkIhNZSmEUjA+9V428J8VeakKGo4dah347TFFJNlQy6Bn/N4m8cbTcYaD
xePvNf0UTQ204iY5nCahgCR4uSC0XfrKIofUibLWCfwEm43gveEDr87yiTOeGr5K
PiVB7Kt1jX1wRII5qVrf4DE4QNSFiNlYQz3+A4TMGVfX+8yXlOFp+JrvqKa+rGlD
nhNHBiG9hpfxWCGyaOkR2pyPMNCLV4/vetJ8FrCkaJ1atPE7XSvpIwVIy99Rr7LY
16wIWAoiH8Vz8TEa5go/QLcEtdxbCnOxBvw8D6FLMg3JF6ln9u4jfk2wg8kqVvw9
s3L2r40EVp/g0DvvNW8gtWHvJTl+AI/cKntqblb4Zdh0R8cd1RD9MRVWXKH3swk7
rZDRAcLzi+r362WHC/8qNeh61rus0OzfZ1WZxOMhGX7Vd2UwQik5a1PDQaGBVcEx
/ErbGZe8KEVdW1Nu8DNT5afIi4mOHcNymWYDvvs1C0yrrcaaryz6EMkxyZ3gfQTx
ZSwQsgV98++FHV4cSBTOrDDLJJa5JZJ5Uk9XND8ZfVz+RqQQq1WQK4zDlfSddW5v
xea+6mIKNV8cKh+2IVjnMtQrFQYUy2ZBlg0Y11uo5gCLiBW2sZoqpYdCh04p7ogQ
ACPkVEHbL9JuLvmhDsNRyDajP10qjfI2UpN6rHNLKLDTXlfyEd4yVzhi2ZpjBHru
KLWo8jBeqtv5aZt8kKs4Ny+3/1hDEzR8fQeuqPMTISf9VMbDBQDERzfXyWFZMlsA
qmGVm4p5eutAKBVlOTR3ADANxBvZmhmHfM+i2vHAIq/WoUvJrFUSfPtqZyd3l7jY
Q5W7w3CmKtz9kvhvSHCevHURlJ5QqnwbEb2YneLD88vYPPVUwdUvwmFh6d8ZeQZP
/reZ2cgXUrmaVfe8P9HioubruyZCU5A8e1LZlB9A+ByyK9F0HbPz2tyBcbAO6MKT
KcVoVXQiz25YNEVpzzclBSPUyWpNH4sud+BpP9OWAPDm3jHjDaspLiVLE8Nrswrd
MWikwpFa2326d1e0chTSCiSvQbskpmhlBUqaFQlzK4/oNFtVNnxFQ7vV1ivKrnDi
1NCxerjnqQEYe/BhWNcPTfJ8t2TbiYMnqe/skmwb31o/hMWq4YRcasfig4tQCrKX
GuYMBsHkUzWPMyhVwWvBm+NHzMGAdw43ssLKCyc99NsfVKnksGiV0fQVkGdDCWdq
C6Vvah96S3TfmG1VVue+Rb2hJK5d0XSaH5VMHpy43Wmf7xrYD8zu0E7uQrwer2BF
pQXkROzLmhzif7+gUkGuHstjReoKesm7YplBAGoLSEi9KXhDDLsNwXE89gkDnI42
wPsVVCrI2rLxRR39QUJSVGSndSiDLmv6NOz/6/VZHXLBdJahKGWI7sje68WFs4tw
e7UDXvq6O8GYfkRBL5KHfGg4DD5ldrYwWnVNYA7ERv5/6dzGNbmI12FJlK30g6V0
25ErPbDkqm99F3XiMdrNYtcyvNxR2d9pTQRLcPrdlBHT4dHjtkBKnLgXvt6vo6Dk
ahUk5ETvk6kToS0/etzKjPCb/k1mnP0T74yWHri3KYLph4i6u1CbbOONnYXi2Gz1
0Mnekh5xcHDLSvy2aP4lHGjOcj7f+QpPldzm7i+98UBcr2Pj57XfJVfcrX2GX6yg
m9VCuEi3fZ4oy77nxJM6UtnMSHT+uWU8r1yqv+Hb0VD7fcFkOeNZWxrmvHK5Pqq+
EPUptfc31Rh97yfLRtbXrcppg2PG7KyVEu5m1w2v0g02l63kbBDxYo6zRKmgBMLz
I3yzURzBwJQMDPjJSDB1s0+9LAK3OsZoLX2OxpFS0fMMURB0SUFBUuGTxi+1D+BM
0rxQIb6RePtf/0U3li1/mIsdV2FPLcMYpAspb1JgvXHrO6+OWEXY94WumOYFEVSt
acLn3l581QEEKlp9Rx2IzCGPCYexZtzy+o8v3rwBd93U2LEV7E5mLpAckPMgAPGM
XTp1X/t9US80y70T7hBkw3JWPcPKHhRzBmR4UNuRmWhjaVnTK0WtUQP1ocnOeEiP
pXEH4GgWB52c9cKwKsa1mY/KrO845Z2MRy11jmVvnCchpS0NVQjWpl9cOHILXQU/
xkq0KfN65CE6/q887iknphJulc6pmb6G3kaXmuxgxFvsft9BpR8MqmJf9wZh22zZ
oaVKxZuxYoEX5Vhjhjc5chrvx72/72bzClyFAlgKVJX8illkY2dyE1qYpEGTBDIb
uqofpQ9qGF/7hseXgy3LlVkALzlYNuRqTze5JcqVTzOGSKvhEYpJRicGB4nibXG0
Pz5VOaHMCOJZIJTuLPUw5N/PlJLMfdokZYGZEnClpOuK+glwTG2f5bhQ0lOBMmLu
M0GNwt5f+2McCkZ5YUiTHNN0VPM7ONrFQWC7ws9ITMuknEqsdXOElj2BCr6wyUp1
h/cR6dzjZCo+FmsBiymTOmR1343WNdntApcw/ic2SwYKk2Dscpd6ukzb5CnGGw7P
0EOl3UhpCfEtvCieKEnzOVhoWDgnta6E1k9pLWFWBMzaKZfkBRgtWiFBzkwh4cqE
d/aFwhSrqRt7BZ52QmUM99GKxVFFpu1apHxR2XuaAG+cpXKTqmAc/w2ys5mU4H6T
QzGN5TszirEEOJMAxWdz/GYrj5MQtApTkqlvU1KCm12jh7ySg60IQA2/ZiyAReQ1
aYHCPvQCIgWaVyD7EOMWreJbvano69vXeneH0ZZ3SmdQqVCYb6A2u0R8eotQU4cH
TSz/B+hDxBPlRKeovgmlRk0zcb8krUU9J8Em9aF0n5OmKQjJSlwbO7lMMRBaPsp3
gwWD98w1btHUBtRVVTGmfL1XlGpMLMto4HFp4Dm0u6Tf8XA1PYMfzlzvnxUXGSlS
3ny9n6ZFlmQhQ8wYv2DgyAb64sO4jIjA742/UUG67u6MVKjYCC2JjzPshPDEyBij
/QSMhjPkjxnf5DCWYtzI+/xQZ/sx9XVRamVA3rwdG/fr5GXFdcDOG4UruiSMKjQE
mJ3czG+gsybPR2mo57LqHV4Fpfz9e8k6lBR5T1HDXUzbkzbjWstk965NMwiQOERn
RMj91XzNQiupbABxyuBrrTk0fObNkJrqYqB7CYSGM8Kh2HVwSvt0Cmt7ni4IBHzs
tyDqMUgH3tksW1cAl18rE2tfx1TcM7tCnISFjYISxWXf45aPW4N22fEVDhUiD3t7
QSVREphStsCbz9tpCHa2rHbc2zd3v973PpDo/fIRApQpx2AhlDUEsBrndzljJUG3
HnEjilupEKTqP3EO8Qg6yy/SJos9g8mzQ8pUsWoKT1i4biL7TjBy+WwelFIJ9EOq
oKOszGnLejmBP3J0YUEdEN9Uz/LNcxxLfGCRJlWS1wJyWCL9ydRST1+pWSorHTdR
oo7YEOj0VMKdbzJ0d4UoO+CTY/i5GtuN/fbHJA9plaDvD9uHpXdB/bQH4iDc9oZH
WGvuolbJXzr3OhCejvTOO+Jv256kmILNBllYcGIhqFWnC6txdFBPZC6AD+vInuTV
pcO3mYJAcMOadIuN3LRP+VfDf/MeKAGKhxMe3xUUfYuJ12K3WlKdfhsDj9TmsCdP
pwRcEISuAwqjGw4udjFNKBzT0hi2ou4CIVHOLHmdvuyxMV0xZxuE99BYY733ZOGk
N5bKveBA5HP0I7FotzFIeM9HleL9YZuz0swYL6pCR5lnUD2TRF9+FNlrN9TjakJR
Jg7K7+V1B6yjPYG3MtnmEpOj/v6+XVJNk4OkUFj6N3HXpJ3ccpboTXAz4D78TMKP
ksPffmcqOPbPeDxnTrU3eU+5QP1RqFaAQqbUmyobdf3DmC2+C9/o5+aQJdHwFlVa
V7GFxw7bYajwVwHcSxSXvqfUG5guvRnEgozmIHY7lsXvNX1/ZPcY6o3l+fOVc9II
tp/unQpLUtiyjnW8EqAabOQZUZBMA5V6lLXTAWmE5B0woJd43gYPhx3TOHIOwrvs
7NtIG5LSSHgMqLevO4VbAAKun/+/h1WhSNKs+Sv/RIbvHw97JiPfxacTxpXADbUQ
h3TqKddvjfytHDkInqQs/ZX1I6UhHiYzDAtP/PwyCTYhKzumtTosTRMQDTQ9CfYQ
RfSHgD6vNzmsr6ISZTaRGv8lS6S86EfICtqkfg5CdJbtW5U9OwRd201cFk9yeRaX
7gsI204In681wdOpgHLVy7pNChEnHXJGLztogIA2NzJo1ZDaSUF42/YVyJxuTGPR
uoSkqD5Ibm3rCdSDvQF7mK7IGuE9VSHljGI4kiTcSUZBvL69Iy/5gf2226lfXwvI
RpgIoORxk56Q8MsVYSQ6X+qlkcecGoz2FCZkmOD/Z2qaKEzZ2hg4cqm3vTqyJPpF
+7ycGdSvXkOxFjY8CZS8/G0VdOZwSLsJ9JI0yT05FR3EWXohynYXf0XIk37Vx18G
7IVcsZ0XQTwS5D33idPVmHtfvsZoHlPmZiwDxuIMiyfZfidl87DrCNcMqditL20+
A2brSY4i7wcR2iLiVCPDZEfEn/rMM6Df0AtbzhNP/zpujJvhSw6NZR6YcPPVUvAf
uuXriZ6pQ66tvB+N1erG/zRrv9YlUQWdc9eunGE2GtxsgqQlZuGvc3Csw5j1hlPt
QptCR7MjPNlGGca1zWPLm+6AEx3PdDUdAmrt6hZ+tCqQmLxHgDT6LbD2IAMLZEZM
zyuMJaoxsIrF5LsGy+H0x6+rFklj72kHqWGrBUCnjVpvuJp1cScwm3uHv+cL9ji+
+3FZRDQMkcr2vvO/L2mdpcmv2St8+WCogJavhy0Ox59dNxVhOq54NK1P+o2dntiJ
UYH+MDMNThM9bGSwMYpYDtZOVJ+jOoaz3a70gWR42DXV6LgWDT70afL/vW2KxtbS
W/Usv+om7f8zXF2Bu+tqpq7yrllil1iwP6duDBQ0g6VOUp+vljTdJEoaQjeXl0y8
lkh0D274x//N9kzBN378XQyVT0i3mKBHCd6z6utzR2v2HvDKc0oGtMvWiK5jgK18
tyH7bBSq+be7r21ftt/tTf/idTV94hYSxErHeFTGIxIIYHxvyirwRkTq1WexPL98
DSgxBal0lyAgNnosKGoSkp+L/rVVhbEoM/NR4Z4OFcyiBkzOFXOcivX33RReLN7s
YRigS+ORV/EPcnDAkc2d8eUG4T8ocVVwM2MASSosLQoWMRsZBvwThXKI4sX/Uh1+
L4Wq6pBzjxDs5e9SLmYNcmr9gmhNvNHyXulZM8CUwOsP0Tb2mufd5jOX6GG20dke
IUcHTnntUGU0rq4KyIAZYesTnOJP8ET0AyS8Lsgf3i6uH1OInITopVH9pJ7WD3CR
m5DnyLAK1Psho75GAEnB3ycl8FA0Qica4iDYV1xgCtAUbFrXg//ILfuKlLi+HLlj
Xy9tFjC6ibfupA7tEA0lnnW3XBzB0jtS8xv2vHMQEGK081O/0EszTSbcbQ0x+kjj
XCRZCuosSdkqc9+hXUcHPYkVMDNlBYXNY9S2gZoUY2azHbS/Vr8IPKWdKgkR/cHE
H+DmEV+OA1XlpTJGW3Jdf8h6VrgNL5GYlFKDktYg91Mke73965o6NJKSvwEYnOLl
JkP+xtVeh7C4YfrFYdpBnpZ1bR51Y3twYJShtnkL/zwNqzhefSGXryz4tne/+2tP
i5ypTzCDMx3REh0TxV4wjaZyY2fIaXJ9JinT0D6/zhvsO1u/kAy5tceyD4p4CXmm
ccNCJiBTRdabacr4+aBzfLIEOnq4dPbokEyWTJFSjbH2f0JHYmYnBN6UWmmbSrWm
QhSBpTRV3VYXts06ib/ob1eOJzadseqsemPC+/ztD5V19o5AhcRp+KZYxmXyASUC
kg0UDX69dzmv5MX3xWZhVl2M7SHTTsH0cfj4ze6c5+4yB7Q6lMr9YaNTC3Fv1kPs
0z17p/U1EuttJdSSJCk/nZ2wh9UPOPegvjMdokpADu6NppSGC7zdh3KzWNvlS9wO
2JkBjmXCJK4PPShSrOXB5Y7KOZM/6N6SOxiOMGI06JoGMnPXi04jUkq9ZMkQqsM9
Hh0587/Vnh8nI2czdwIEVQ68XmyfKB9oXKNnlu5dUQJTq6CAOKcIKT5hvwty9GQA
i5cwcSMJ5iaqOur8mOyzcvwbdA2WRt6ej1sfgNLVR7pdzlmvzvIzR+NK2dLOAlfq
g9Kf5QiWC19Y0JOp8mNL4gR5ekttVhpBwEN0d2UlqSXsnDXhlPGaRUugW76uJdSP
Mjo1P631MOzLdaEomMLmF8THv3q+TqJuZvli5NGwiji1/v//tGdejhLPAvtjZ8Rw
O1DPrsjFBAojM3X8j6dlrTJ9GCTBgUMJCHEkGa+Rjq5grN4QFIYWEPf7v2K37kF0
ZRFJdiF61TUsTH0Ck6BSzC3UoRk3Heo/c1qxV1hE+O9qyu/1rS9xxd+/AQfZQuGG
iyb2WbA0GxZJbwcrjtj0BCsyeH6xMhjRvCKIwWjjrRsrP2V/c3p+uQZBLP2Cmx7b
deNJvha6VPGaARHoMr+6QhwFfVXf1AS8UVVcHWaSqPm85jvUgqbygntvY+0xVdj4
K+KQ4CAkChu2+GdMX4CjtRknYlkZZn6ZPxvqdTeYZO9/IDqjxyDNhDAy6OuxAJHa
rt7LXEHU/0Caygpk8yyh3OtR8Y4jexKjYWJfEeMFxV2RerVXLBLsFVKqkimDaE6h
lETYOCVjg0KTHQCJosi6+FBMYrBBtZ3RDgd6iMYL/JZQJcx6skOwNMoi6I+7gBJ/
MsMdXXuowS+j87DcqEwARW1qEj8KOzwuHMUeDy3eUB7lZzi+YnLqcbEOUzQK0cPv
QSTp+JdOLQxKWenZF9y8iYlQYUiO7qqZj/+XibxvgwO7NELWFLNehSHlzbSRgQaS
9tDs8EenUuSja24Z1rtZF6csZ2ssP36ozvVRGquTwCF8sc1V2edRYMhzCeK7EuGm
2NzQA8I4WpdkBpgpUXFX1BqrSrLOgfbWEtzCElAUNY9CEUDqmJZJ5CQskYvqtaGm
hBufFF2RpueDPW+LxdLZ8DcPlshf9yPYvitAIazih+1u4yns2VEOaduwPeW5kEbc
slJ2hNFyXvc3+fbsl3gHlvx/Z8m/STHewXSZ3QWVBcpCa5a4XhbfI7YiVO9McfIV
LfiH7LwIEp38O9RK4fsZpPNk1fKkgjTE0MxSDLYSfPQGRoR3ZYFGQ/GfctqY1JqR
pCDt7Kw8CHdgHv8vR/b1+kejDkSbVYigMx4qPdfeL9JkEEEGKTx7saRw324rOdR5
xxA2dyThi7VxTOMm02GeeQWr/76QmOqEv8pimS+b93PibirIBgA3LIHY71x2r3sg
s7Rxnlx0Dukzr4KwpjOjBVmONx3g+Pn96XM6pjqe9GmYco/htB8cqQxTSPS0BsW6
q0kMkiV7FE4HFhBwBd9AzjR9ysLizWWFhGlUcDdG8YcL4741JIEIyYImNZLdGdiq
SRItR9MiD66vbX639jovJ8zNkizjXwW/XfOb9Utaw5fwwULNg9l48qqNOT8gvJ3V
i3ybdqb8+LNT7tGxmuE0tL13rzDqd3wT7pKTFJGJIQHOYBMveKDTpRZQi6n6h3R6
BWWlyqpp/qqD04PFIxWoZbQhHPpKbubRMlkvoWDDRNli+0CnKJosWfRQgqqJTYjM
nlRUw98ZTBtoaC/JZqKjs4Pehls4SC2ykOe6llNZVSVF99e6/rs39mcdInr9renI
0zxI/AG2ueRABLIh9FxBv7kFRtMeSPZDdhI2EwV5uIHdNbonnyN8jfJ/6b2S0cgE
VnRSowUZb5e4ne5CajHj/hJFunrihSPKzqKxMA1QG9be0UG2OPMKqwfrrwOnCYy7
N9IcoZlUbQ8XaLjkLat77g21nyTW2VrllUtYYulDR4i764if1K86A5fpOfV1R4Xr
71pTjcnpwXcHQICgPo1/LeN/aZwZXulRajOzSu7EkwursdiWcbTpHIanPZO6kdKS
/SLAJhjyGgKxfzHzptlAw9vSb1/5GnTci+FHFQNbc6IR044E02t02vjN7b77NpDu
yWH+IcM+AYL4JQbIgm47blCDMaBmT6LpOCFFbM078tT9sqRGXnPGQXrttS1na/lq
WtejA5KjUVNaKUT8/j+OF78ewAVMJ8zBDS+HFxwfQzxuTVNTP7prCmbbg1mbpJK+
Tb+ug26up+grJaf5jl5OZaJiVRjINSAnqiyBgLkFSJp1NtdVNma7Nl+YrQAuVTRS
x3bSskThdyXJu3an7eZkwPHaFdzAAPWv7Pwe93JUZkui+/qMSLeLH8Jmb/1k3Snw
lGC47Dbf3Slhnp39CXVWiW7vScHcGE15DKtWNPP561kwI8xWaYOyqZ2sSvCnhasW
ZSy4s+qe4KV7JpOk6qpcT/vZVJL/xqAluMV4l6LbxlrbSO8uCsr7xrUwZVnW3Hxt
KjU0fqny+6NF3D/dcOnIXatbcvzmkf222FJFxTJgZsYPh5InnKW93HLZ6EHClJkn
lA/dqNGX02JOe5RWR1hSk/HYJ19yjUk2A4i5fSBPz7ybuyZmsifoBS7f2zhImVPS
ljvsh+MEMtL2aj8BRKJUQIsuo172eo0rYnNy4FDSpOCtu638xrREjdRGravHtj5B
x+fsRtg/CjCfuBFcj6hYAsP+6rGQXkeHMxYPwEJVQ/rHobKf7jO/3cC6Y6mrPwvL
H9Ubv5/uEO3coFRanLKekjquJaVDbtiDq3WBgXuRgE1BCueGcvjeke32ghXNOm/a
o2CHSKcPECgssvgtcIvMnT0QvAmn5VeG0wRQd5WYsG8LxYcj0aDfiOK1bjraFCE7
1Y0clksABYs2F5a1pceKvZ0R94ZWjwqBp4tOKTJaOLu+6D0kVNVUM7n1gd0KO0tm
M1Pm5AavjGOiGrbjsh+EIs02zUlH4DvhGzUYAmUa30Euyf0C3PrtpWX/UYDXrybz
C0UG65hVUveGWTfZr4063EHT2yxfYxGfdvuGzVpHgHzt6BY3ccrEdjBFZGB8YzOe
LAPnYaiMXu/eSXrgiXxYBiqfzj2iwmFPH+DNrxdTfeZCTkH9yKQKN/uADSHaVN3e
Ino8JoEp169wDliww7RiLXyVCQgbFuLP+Bjyx9483H0sQvTKqG6PESAiNecc2G+Z
6Sb6ynSGbZ7jyQUgEDfmckNLvXmDYa4gU6jmNabix/26QORDlkya3enaeK6PVRwq
i10zblfK/d6B/xL18qO9ekrkNFe4yk1Z8+3oJ1UzpprtayTW1GX3aCjjB4GKNw4q
eO7yGX26Gt0H/LhxjZ3z7jmoCmYFlqg1HT081R+bgNQtmjGUhLMeQXGt+xZEX2/O
eJS2JW4tVoaiApZMQkLIRhu81uC8SefogCautR+6agJSDmcWRQq9l3lDshCBPggX
eQtFDM9e/0ST4s4XLCn+DJZWg7QG8YFUe5YHUbXT+X8MshprYZDl6jv82lfR1TqF
l/ngRHxOjd5ka7pAX4OtJnYJHoplvUmHBj+zwhRuybO10lXifLoCa3e8/NIyCqMt
tY5beZDQh9rYiyJWDbQadOIVxi4qDujwfoo+7m+a3E4F2WGnzM6C+3p9xQxzj9av
ytCuSTQb6qXMe+x4j3FaGzuqSz3lWQafA0qWDDD6CP2t8ALdqd/4iuQdkTbDdvte
J4WvJuklG/jD4Y9KXvpDjQpL8MQyJvu8VhJ8gR+JqAk6sHDfDuVI3lremgaxU9AV
HuCWSrGbjwgmEAR0uPry6MlbQWCRyIozS6q7Up1JeR/Lzso94BkAvRKyIddc/Xxr
+ss2ZN3DqyIraXtQjjYtz0s+pe6g3u1oELxIBqCLJ/R5BwKXrscpd+DZkaEFpS1i
tlVOX/VwHbUKDKXB1qMvOTk+ySdBc+wMCryzhXTUd8s3+dXQVU6aJXPTYv1SSO17
oqkUMAtZ8d4liqOKUpDz/iYeoETp2pCLfsdF9QlOgIE1rK4K1CLmOdT/qyxI7ou3
qJv4N/hZmcRSNYgXtKqkLfJ/SZuyHBJFrzsVJgg8TYzDyKLN5OqjBqh5GNhiBgBx
tlJD2zGP75HudVDUBM4Ixl67QjnkXFDg184v7GLDjwJ9dP4olG2VeZ0WbXXg3atZ
XAPywESXKWQIPYvPuYgk94aRosCRjTYhpOzywTYxvVy80V7yIw2Q0u9W6dgnINpz
0TCbMe+06QgTNNwzJ39bGPsKfYAxKnscnXI4ne8r7OElfVdXZPevzVixixbbgnms
hOfwkiDwYrhWLPFY/6NUVS5FfdDEv0vNCRJytvME2h1CVuPq54ML9CsAem8GF9fc
R1ESLAwE/J3c4+78tZ31lovfPpiPnONVqJ9m1gIeGFpZEvMQGGSSogEnEkuEagj7
Q3C9Ls5uuT02FSOs/xoGhxuRnOp23/xFOBkCQs2y5ajx2VdnshTltMA5WJQ0S7Ky
eDFW00z2ARKK9rXhjF+FxyRtwkEAEriUt8jLKbLisgQJxKpiD5oM2RFPKSjxBD7u
6bfT2pkZC0rALKJHVQTe/QPpxoKTiAlYT3bBKmEfE9g47Ddi6a5N6UFKY02RPe7r
dlnNcKs2H9O8IG5+JFuoJHgtfi6K+DRu1a07CoWBF5e/nnE4TYGGQ2zDjqIGYaAI
AVZ1KHmpt3TR0YoM3MOd7WYRZCpLoxhP55VwNyXjoWs+b3XnLQoGeK7J+VoNhaGx
1Chq8QMXSCcY6eBXHkN/ltg14/qumkMdKBUVqvBk55Mrm0r52eF8LXCwc7+JwTok
QqP7QiV2h220mDaEYih6eSywk41OCPgP8/Ss1GmjQgFC20qdNYhba1gkb43+iTKc
Et4yBnD/pzZqz5EJwkP+vVuEM9YEgIAoQZLN7c3lR/ti/5AmVy9ddbhWQFrCDSrB
lo810aYVtVjWxr7HbpUEiyV/kCNHMhyFGV59ftaNUNTJJIJ2Udj+KTqo2g+1N4AZ
r0AOjTubiptAedeGWOL6KlWv/+v5FhQRzIX+Ixf21kWj3sEWhba5YLcxMM26gEb9
p0egC59HgXacghS40Xd1LzbDUJYtbgH6/3l2JQOzkVpYCfOYecEsoJmca1Nqc267
8QGbQlCm7DQmqvg/cBxl8S0THZqEOH6Km6uvQCBshRRFTNiNsPRRy05Mxp5HT057
cM/0fPwNjvSq5AXtnDDUQSC2U3sUumW/jeiNeeE2QJEmUs70Iwz0g76td2sUyBV/
YnwRlqv35AQpRuaeEFemMu35SZK4bmnEVjZnQlLx//JhSWNQkJEubmSvRjJKLxwE
fC/BfxYnyoC86A/chc55GbZ9zANAM2vQsg9xuKrMM4GdGWCnFbPXsTy+rT3h2edf
sjLnnBdMH2ZtI8CBAD9+1/53p/oMYnwjMrDBhiYrY/uyATR8bga3UvA6JuGqU1bV
CbW5HvR83429AWNnbKFTeSjb82xfA8WpeI9gzyKgfEPIJVYO8YYStlBBAFDoQo4U
Jewg1sqTu5h/4QB8Xgo0abbp3tYYLUzskboVGyIjoJlZmfzIR/7mz7C5dT9lNC06
MI+4UAuFr2kc5OwFNQYdLay2mQG/AGydLKrHk0+VG0SVh6A0Mo5jqRu5aeKGOCsh
v0zjYFumrqN+anvU524jKyoAVbS0UseRJIMXT3Vdr3F2QkHDhkhbMIyJilAjnExx
6f34X1/NAzCrfOMa5kEawmg5YoKthm7rxB6w02ed8yw+Rr84jyw8ie4ZdJEC8F7P
qaL4bJyg/5TdLWkdNOyUfg7wF71Bq1kE+kEBEYyuPimL3g999EwW0fDtqYlCNeCd
as+foLNa9pgtEn4PJvXzGYk0wV35TheGLvT0XFP4o6lVR+WKClXFBP7fBxI+0o4f
LBoDhi3lbfgihtcZaNYwWDpGZqq1zWUuHmJRgOosmbK+PTIX10ty9jiq3utH/O+q
jmCfy0diISWbKFSITvYyzuGn9SQb5MlFQ5lwpRL/kGq9ELOLxbXFqTYFzHvkdYQ2
KBq2nYE1Ms7JTSM1v+BL37aawdA1wQZ0siA/Bc7YHLmuW0hqvZFDP/F8AwOC6Lrq
OfK+jBzgKpoTsKKMXowujYgZHaLYN4FQnP+dhLmIvQOqMDom/+BoUyxrerbIBnzD
jI9ydzOzJYgQ5S7Xhz8xvwXhAThBOuzvxb5bGz/hqk/K06c3JHMNfeANlnRbvl5S
FBymxCHbD8hCWgIAsdG/+9w9Yv9CSunZs1KBQJZlHaiib+h0/WOZuIPpUkqKful+
hnSrttLnT6VgkcnY1kPr0fyfEzjDrw7qqzzytEcgHEdWVQQfEProKJxpmMwzDvdu
neguvfEECpCmdPCuMNeCDo1hweCfH9eOez5VTTDdFQvDtJcD0BWzWrrtpF20Om9d
zFBy6CbadArnuUxDvUnteO31V3lsK2w0nD+XGtF4B2smuP/OPNrwkkHFNZaKHs1H
uUCpqayzpdgqH+zw9C9HbkLgLwhRQ1OJD1WUPMo46ApfdcPhszvPLsxbqQpCY0Dc
JbtYgx3kGMl9li4YWaqpmyCn+A/qQYEH+9AJFiXy1wb8AJ8IgMZ+DTfz7+EiPqBi
nf0F7S/kUG5TlfURE41PR6kefMW9saKzDxCjjjiKbeKedYSLw0/svaKI7lOjstui
m+Q6jYmovES1vyk0fXZTi2OF5brlYGkquroBdvhCkvFdMMNi+3t6kDMPnHSUJneq
xxneVIGVAuhjMAij8x/yP+dFAT8dk2Ia3KMDeQieIzmZtiav4nt22WDnAkyUvXt4
zwIa0EQWB8+YMRnlT+HNcGqaER4iJ0vz7iRXZsdpZiJz+aS/f/lrYQET3E2hHukY
c67P/JH8fNrLX7weyqvPqQgaCMfXT/HOMDO66UPwQUoSOa2U9GHdr0IiyPpG3yS9
arLLlviAp+U6zqEWqXkz6xD/b/pHQlvzmT+Iw4zK+GCx8rJjOWV3qPACH3KxtA+g
Qzl0lzYb5Vf1a5hsunkhGwQTpFeRUDIEh1QtbilzSSsk4KGnGrV6miiNNpTfQyJ0
kbhJtM7heiQ/9RHhH8Houh/Z6j87aCxGB9WIPsfwcZRtuyM/Hw1+Nom/Yk+WmslS
NmL8wZMsmt2jCD9N+jWynS0Hnj63XYMTPe1SuuNpaTEc2oj9XYaTT7uBXsqpol0B
Q4LmNGtHwRw6J58PGEG7zYZ41X8fV/MDPP7q+0flhAHlXoYOtuzq2MKT1EfRiJuS
RKwna4NbxvLpP7QdwVLiJClt9bpxrAGQVr/V/jod/AXlB7ZSZE6QGuDYSMkADXY3
Wjf9g+n4k4nsn47/9qwyw/Lk48RBouJ4+6VWS2gWIBvkOhHibS/fJLp64QIgsnH6
gQ8VQN9Ec5EMw0qRbwhYT1sg0czxN4hAaYjkwwgBJbKoMLBO5vuBSjs6iSAEicR9
0ra9TUM0iwGn9YuC/edPD+PpXzH4XhUItkdxqb9l9rZ/Qh4Z1NeRCqIMROrRlGHo
GHdA1RHNu433oAduRfnHFBmW3wDt95yO2iFKO4PUNS2B9DP7d+GfuW3sTF1KSgv3
22/PTeUsZQVG32bs3aSnERqCLh0oczv0m7mSbNeQbpb98rfxEuBPcd+D6/yWjAed
m+eJwjfn9uai5VmURc97waL9Iijj4H5xG2VcNkNAOQ1DVEO7rQqwh/HCMc3I2J2R
5QvulpmU/NMIRho/o3PpDEVM8+VNcLvx8NQ/vyWAtDaOHur0joTDPaPrbLTaTicI
Ats+/VENXQ5ThBFFVJURCaCuLe3ebx6vqYqZ5pwro9Wqh2aUFB7qzSMf0RXaeTLh
anqVUj9tbtDenVjTIjsvd+AwTLwFnxuyVrKoBWLS9gkxqqJwU1IPg2o+laWc7pwq
acPQx/u9LTf4uY/BWBkfPXQjGLOgkZmuhmEGAjre97yf+009Y08UBLfPrrhdYBF2
QkOXS+SE9Y9sZdKVaZ8OJ3rfr9/+sRvSSqVySwqxl3ITwr20w0vWQIkWVd+qG4C3
9UWld29qJng7mv9+gTt9xbyojoFYs8doe3oZega3e4gwohoqDGmzmVaeMoG8R4G+
lDiENEHH2i8Oi6upfqSARBY806SaAUonyVNcGUmaPacCnanIv1yajIcrsD5RF+Ah
YAYj95DBvQQEE0vtBAltncDIPNH3/5v2uttmeyA1BcD1MXS5T2qkG0SeCvarblQ6
4PhkjsJkzlkxgbZfqwcsEpP+4LM7ke6DWNfWp0URznY3zO8sVO3ITNqEXUKh2sUP
dbip7hMo6X3cdekeEBlMtBFwIp+YZEdTJnHJjP7SUP3YVTUnAoDrYMaylwqITTWo
tvVxORUNmhQCidbxE7WPjfoIiGPCylVR2NgWTNUBX0N7nVI51Gt70zwtDnGImT7+
fVfrD8SeJiSGnR+DR2cWCjkX8R/sAGST7nlXYebPz0snbUYPo5Kc3lNJd/P2gEGE
8CHW2RieIUCd266AlvQMvNP13Ei1qw1Jo50j9tjeHEngn/4jJuI/twXgS0hWBCJd
cmJJ+vZUyxTf2fKS58lXg7VpQFtMPWuRkHZgwIOiFbPGJtHoHLfZB5Vme4ed0Kfg
SkCpnoq5Yb2DQvgnHrTiq8E7mG8Pz6US/D5dmlSUoZuBtMfHlwqx7ZK48mU6zWy2
fnI27uG4EKJvFEK+myera6C5/XJ2TAHo/Z8bFL7xbbozQGvNnXMrW0VEMygtpBR0
fsFAtdH+GENLcvMazFlmgz7J3jCnG/RpLKlUSd02vRfEhRJwruCE8VbQZlPle9H+
IRogtSiJCZMzFB3ulAiPzRzEuLQdYXM+hPpXkcWVWhot5hz1/de4We1ksbSpmGUD
2rSSEfg8SzZl3Fk71Fy2/1O3tTE6DFZ+5MnOpBa4okQgPyy70gGU/URBbQFLrjQJ
KlegA5+eV5jnbNFnB3BE/+ojAmkSx9S6aGcYbRaWACsR3Zmn9zcHdD+OvZR2kCCN
Jnosty6XwPt7KusFhxTXfKvlqGnYXoDYuNhKmw740/kJoivKvQwWYl38cuwJBonV
USUyGgZPBOPXCLMVdoFYIXNmwFqt4WH2IBQc1AIcNOJW9SQ/olx7X9RAnx7YpIV8
lAfA3y/HdEqI0+rUfitjoiyky9FJoxTKfOrnNQYpLn9uhWjUJxWQhcZuQ+S2vTjj
8g+YXCJ4dboPnqvGMPP2nYqNbKt+Asd9Y+gDLZC8w6PXOLfXSuZ2z3fpy/Hy+e7q
fMVocp4itrsfpn1m4SSO1MwjcPm65QN5XRLOdVjvIFd5tGmVH4C/aZ4Mo5nPNlGT
ZpjDLI7Hj7OEUvZwrATOgCI3Ho5lcx21zcqnPNjOnOduzHmFHnKP7ZJLVUM019pK
aFIJ0eegfepqXhzVewqB7/LtAaOazuoG6oaP7xHTzb4BOW0zYGyK/USDywsq53bn
o1YT+kq4UlR5gYJFBoE6FzWASCxwHopmpxGfITqthjGjHBl+YvC5kW5NY8kxrcfg
vH/KXN+CJ8TJqMR1vklpaD/tKzk75IuxrYAozjHGlnbcrSqSWJ3cZhHp5w9b3kV4
+9vaTUkwY+kHnqs8AqG+34e94T8UCgZwl/uRKutIwn1AeRuRwZ90MQATMgtDNhzF
q0WLsXF3cPlXBUmjlY2kP2frxJnx1TuxksC66Asw7KtHxRAzmbZjiuSTQ67LEWGw
6LZQe/zZbo0QHuhTwm5rHGxGM146cx4J7gGoRDfj/DED4pPojRJZtZ2xayWVONAt
iIcigt451faqSU8sWwQCiJM3iKUWnA9NGfNujX+i7GrP1J0H9L2pu4xFjImMC2iA
16R/EouPW44RcCg9RY06taLu6J2cdbnXWXBIFcpjn6XJpOLaUQM3Z3ACG02wqYUg
uelRooQ/lcmlD5+FjC7/Xfy2tdseKQA2i0rzDZw7+JTovGrIGPx0iY/xb8CcjCxz
UNCnBhlVA8LQSDAHykaZ7CtQSgkhaKamWRv5MAVog4BXNgD1NjHdIN4E8fklVWVA
vNWyaNbTDTXfIE+fAWc3jCuRzejPtcMTnf/bMTg0WTq8k25HZjqO4CrZuEjI62ar
sCH9FXnNDVq6ql3KHkbYCGjWXSuoW0Z3LlFSYIzWGdHKq/JH5X2SRcLIASoe0YkV
2YQNY0V12cteCrzZUnhjZU/DolQT0zo+tgCQPRdDuNVolwDU6n2/5KGVTX3JOY6/
xe2poFkWFT0O5W8uQBKia7HH3uEb7Gl28MTP7vDJotTC3eeHpPmDxT5mWdr75DPX
da6gYOa6q4lm82aOAIhRAo3grTTVL4wsC9VgKuCN7whnZCfJOkarV5nleRpxGRDl
HhTZX/C4c92CJTCl4pXI0HStE7RFWk7kTKs37flZtlAQWz+XjoBhr8v6rzZ5rtVW
Uazx238FmDYOxbo/PM8PrhGks04qXN60vyiIOUuWn2XgRJ320w9IEN7V4vo2zUXo
YllkDeuEgsaInWqVNgrPkvXwUw/aJ0mWjN6Oui9VuGnOHc5dAWHO9gezi1p0D2we
279swmN3USUc/zlzxUXs54/CE98Qa1iwnVH3Wvd+TFpTWnufcghDn0Sc/H6BzIV/
/HY1K2Ceh+SPbxhyprMmmA/62XYfjATM4W/km9QcSVaTdzJqI/X5kuXoDb8P2Jww
AF5ythyIa9EJkme+DFCrHDyOnSAvQ8bhTSSE3Kcv3HjdslmPfe2PP+ZhA9vLTYqi
MAPJJkhFyv09C9VZgi1RKIrkIm8nXoPZ9b5RKL9ba67XftKAgjwsasAVQFGuGKZs
iE89szSaqDux6hjY++SVuoe5yCiI2/XS50ujaZqXfCuinxNmQaW/aey/3c+A3mjt
PEM5o5oJDCaJDnA7FZJY+pocJJU9MslawePuaPnp/cLM82kERRoxiDCJEWOuZCfG
1Lt2sQP7DlgG7/lwG+aoajFUY/row2Pr8j7vFUUHRJhn5yp2daSKw0zQ6INM6ieU
/PnsKws/+ZS+GA30fYycjH1b/o5h6feW35jkzLMjLGtEM0GxCyx/CLXlkDpMXsZi
5VhGuHb4F6lrlkiuKbibfA==
`protect END_PROTECTED
