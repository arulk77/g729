`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqpc6qJnRUjYzv/nz+ykNGDrwOotnJLIVINim/Hx2smFe
oRgFkqgjY63ISLfo97rWwInvPGcR2vGUxesjlwh9Co2f1EYZ0BuJyo+4ZlVxEQ06
/5audBOdVmUyMQSjlUp/phQQ/f9ZpxT+kqqulfgBgmxBKq4/fzJhp/icCR6J0qgu
jpuJSyz7mfwBwr5yy0vyIc0KB49u77q6qjeYXBWv9BrGgJwn9to56aiyQg3ncttZ
zhwNNJfIXpKIb4ZoRHC58aU2SBCIxvWY+pcyl2YvJ40mxDDw3oKqX4XQzkcBY+Qy
SHMXci8K4AhVJ20q1svX7mBQwc40UafeuHIPyujqfxgrlnCATZZmHUE9XE97qnzC
+/yKaNB0UhGUg5mXrnplfFgdsKcuUlSCkcgiPjBLLEU=
`protect END_PROTECTED
