`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJnjc35BOt8DO3dEOnVmxTA7UplG8VdPrZCls6a2hv/U
eB+DYwaaiDDfy5rKtfpeHnS7cVZpBS3SuXQ7ln99/Wyv+dNM4a1e+CS2jU9MyW9z
VGvB59hp42X6G135a4TKQ0GMzqidiX0JEbgONmzJALpk+K5qKWDUpvrMrgNk7y58
zcfbGjOQI9RJmruLtkZugYkWNPAf+XRN/fI8vCvnuosTRp25fHHgvocDBF9m4JJw
`protect END_PROTECTED
