`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
av5LoUX8r2zQa5wkcbU7hH4wKooeLFRbKDIkq0qyumsz90VhqtdR31j68sV6L3/j
LRLuApb5q/OlC0wQb1kT0apEW0ycdffycjMGyVmaSEbvkFjvZYsZLiVt8EpewPqQ
58Hol1O4JNdxqD+C6tiamLqrKSvlg+VgEB1y8OyfWPeQUa3/tA6cMNdzCpaUOyqk
Nv7x8wWEQZ32F3ED4D9n6/r0qY0vn7JP5ANDPW7Ee70a2ZbE2xFhxmc8RgiFUqjS
bhVGS7mDHAMTCHpw5rlyrUBJAEpLQ1+e9+JV3sFYHLD8xy6PIXgSCFbCOgNdwTgs
sRGQDQxRBZuNCeYRJDZ0lN9SsiCKa5iszFLFVrioCwTe+DNtjsVOV64sADQmbi9c
JDrAVA+Um4jVkL56zu1lXR/Wgnq9vtp7y1/PRsme89OwmjbPDD2LHjiYK/1G+Qi8
b1v1HL4lUfj9SZkPFPmOzA==
`protect END_PROTECTED
