`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ypt+YGyT02GtzUmmtyiuG/ydLp/au1CUc8uXLAKXwRd
T6h0qKWStvHg7VgFuHRthG3pvv5XHz+tTlpMhsTKE7ocErZ8igJXYlGO3tRxA5Mm
DwrDzEf0WAR3pf4CYnzDssSU4s46UcYhvTnwp9DE2XxlEuW1c98cQQx+qCnX0xQB
My/EHBzhm6KtNO42dM9UiBGydP9PQ9go3SIIRDmz9da/PdPewSGOY8ejwf57/j2r
i7XdSGafnNDFTn+PL6mpIfYo+m8OEJsrw7WT430m73ufptN2qbKGj6vDBrdjAgEj
axMotKGbHXsP3HIFrKjWjlQC3E/8aSDZx0M/xO4Qlwv6s4v6ccdkdiQfXiEaxNtc
LX0w72pMhUja5ptyidQ0HMvXtrQtPFLfHoUKZOSOQDm4RupbdrC5WyI4uRzLoXKz
cACHpRNWS6RF0C0cN7zOaigHRcZBFRppgzMFfe2e0aNnW9gwpsIBOyHAC30VG2kS
Xiwui61y9SPJZ6Mj4hb+CEO8AbSiU47LF7xIEzEE8ZhqpMiBNlofKLqCiJEH6Zjo
3mptPpwQWkTpdNwwk9KQ1dQmJIhj+Z9EUX1FxvbOTumXbX4Rq0wsfgVSM37h10iS
`protect END_PROTECTED
