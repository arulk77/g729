`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePzyFVCab/RsWl8FFY1+H2X3vSqw0c1DZ54UpQvKD4+l
cDpH4k6WD6RPzq23EVSZ2qlpHSUH+F8nBxn3BISYE1E2yzNIhdS838+DEyi01+t2
iHq0kau+15qdM6eIcCO4gvl275ynF2WleFd8KSMDLme2cdCkIYYdMFA1SZpWro3W
U/oqr7HyyvGjYWLZ5OfYKuwEyGhCnJ6RRmWIUOJq/PZBDnauJ5MhgYkS+B9pYF3r
`protect END_PROTECTED
