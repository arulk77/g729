`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Nw2iny9YWWxbi2/rsVQfOSmxj2foZv8o6mj9vFqrDaxo8PIf+yQiV8ebozONCOja
CKZsGiBL7i/uzZtx6pKGU7oE9oRP/cTOXP7ujpP+HtNzzOuIPUzVQapuWv2ZJrMK
b+90xWW0qkwqkejuaFf500qRv61E6sgTRj4v2QG6sPXKf2X/CCQaZvNrreTTawuA
`protect END_PROTECTED
