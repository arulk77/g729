`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4w5NRSK85txeU4cXFnaoVqkV11m83sK9b4e7rAlDiMAk
SazDhsZwQqqRtCW9s9TcrwPH/h//4TxO2rwVjT+/LUZZeJ0s9KsiGHWqybENJvZr
h2jWr1kE6ghdisbm416yV7Y1iCYssq92KUAJ3jZstfFkDgL+Xzhk8qY41hTH7TLg
9eogVI2SBK3/RlzHdPWHpSUt4I2kOBdMIUb/BXAmWwJUJHE9nN4cg1XPe4usy1m1
M1jSfkbDkQDgB0Oa+p7+vmv5xUk/iHaN/eIXEklC9tFHrJlFwsoM4nykxvxIOYtM
lYCf5T6iX0bzetek23BcXA==
`protect END_PROTECTED
