`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBo0Ssfm2fD750NFi+f9PdiOio1e4Apu7hfqgc7NtiLt
O813J8UcW9vySBdUhY2EwIYIvlyofzvbJ0yQE0IT98hVjsMkbiFLrCAZsNAr8/Y1
UmtxISpdc0XgPGBBZUl0wIDXDuL5vwk8eK7lMYqANYCbrTPxIJxyxbhiO102E/mz
yafbXLWMhkz6YejOeE75yapJF4+HUbgZ2f8DRopLWXYYvrL3JWrfLE78hZ3YPbli
/8VNyIqqRAuIf4/+UUYsDhjxfCpp6tkb/11+FE0uRuj4QsNLIYyt0LPhoBV8T8EH
daSlsgr+lJWwwqhbL7NoFg==
`protect END_PROTECTED
