`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IoaQEtWnqhZxsMC9miFItiExDBQKwZZU1YaL0AmkGAgPEslkwqk6kJlT0js4rHRF
LpMOWWqwpPRHJfKWRqGX37OnlypWrbxLzXeistJ9md9f/pM7+dz1oqv7OroDRMJE
GoWbvRpqyDK0i0AujN9tmAxzsouNZ4fhiw/8/o14shwuF7X1sHMuhVXN3Xzeiyq/
UWHuHeU0w3TD93kSz71d0Ef4kd7bivuMXmg7jl0lOdk=
`protect END_PROTECTED
