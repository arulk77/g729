`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNEpGJqf03RN8EgvMg4eGZ4hK3271USmC0Ve/QItTiG9
gOVw08kQB4Xpunuh/SLfU2GszPuCDc5MwF2Li8kwXK3QOFW7JifM1lorvCG2CqTX
qLubs6xUOnqK8k69MCdhQ0SXS5OiztkLkWiL2pEMiwGAF0Sk/cGhjMcxyeMKjHwe
miITv650FD0NCzRF0R3jJEaDFJBsopX13iXMsiZvQm9U+TRWd5UlqQsc3PauayWe
wHZzLEOc4Sb/0ExwH6UBuCcvnq97MVyOVJQlfE4jQYE9sFo4zW5v+2/2IWZuTT0B
MCUGSg8F5Y71KknH+dMUak0H11GiLX1+hZxUqLvWgF+FRg+Ffcke2Mesc9a1yGUG
`protect END_PROTECTED
