`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu410f7LdmsA7vemHCs2TewH+57Z+ogE1I3yJ+K7eI6E8Q
jzMcFIazfPi2BPLBVKhxUmzMXyYWkUhQE/AEPRzLQKaagXZ7rTSc497BZCw7+6uv
Z4M6Fq4n0bC50q6LHzge3fLcZVn7ENk0I1axNJxaQXfRE17+lRMNWh+8x1DKQdSg
CmZWIDDl7mtBY8a8Yj6Y2PqsPrDchrEn0yh46ahLahI=
`protect END_PROTECTED
