`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFTTYixzewDAYXN8X89osVzv01WAUz5UQS+xchPtXO8q
RMs6MdkbnK7jqGM/T+zYSSdwNsF6PxkNG+GUrQqAnESAlIiZnEH7iYBHwJHAOD/x
q82OGkHULfm2HHI4JAOhrGGWro34D9Ih87o/Ac34h38nJK4+CsTLRRO3b+GVYbwb
My//r31d5Bk+0FWsqmI8TWMB/jH66d+St8YC1UUII5c86bPsREUVg9MQac5u5RRO
`protect END_PROTECTED
