`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vYAyRVA678lidnrpxgf9/a1SXRW2DyfSyekubV9k//ce0EZ+dBZ9jmf3N6gO/Wc2
fTQCi0vTTlO7pLwJfCZnoDdiaIz7cHWkMx93N6CasUweMiZsmTA7YXgwXvv0x8iz
fefBuErEjvamqdWIoUWcTGw0MM60qvS+R6t2P41Eijv+neWt2r/AZOyiXncuLdJr
UfwFBLoLxafdID9mHku12K3xwrijgM78A8AgvDhTojzGw41dOPvUAX4ZtrvfNo9J
2ufVPQlzVlsTczvoOQqwx8npioPxcg/UyRBnGrWwPrg5HfbhT8OX4SO7upSMvYk5
BXPsPHozeMBmdQcI+4AiIpeUEWPnVkWyrDnAWwqzrEA=
`protect END_PROTECTED
