`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xYa2J5pldJ+QMZsHPppw7kBRpUAiQRRsFiGbNnN9rQ+JOex8/68OX1YsRnmh/G+I
zoMOb6JCANtc+ii4f4zbD++yvsm0qTmVvliJZ96Q6OY0VYwIpUIemVhGdSf2Zycp
RoHUSWCeHuwj+B0x06/SRDnuk20aqlZ/WqvmiBgwjJtl3O09zscwnV+IXboePaeH
sbwJJPSdtwstTRZ6NKQCDj0WluqsxMnUd5NRROXKcIXOyDDrwJ+1V9dxjWcvTd6k
ujVmDeDJDVgFTLaM+ClrVVz4lkvjkbjjFh7k/5gAs0rM0XCIU2jxF34w0cfOn0NU
j7U192xKy1iLlxlBUCO4WPmH9hhL64gcgVG4eES42jhoYIIbEw5nZkTpfvGX0Iw2
`protect END_PROTECTED
