`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73Cyo9MnHc6aDVxmgiUZuiy9+lBJrtMKmG27ki6vHMkgYC
7HW3fTFCZu9+Q09SNGqRQtmPp73Y/tiGg8cNMnw2LWdg8ZauiKqo1N97xJm+Bpcq
1Jg8oA7+vNxBkGzP5ym3djOhPNtpaBtCjGpjKf6L1IcwWzMSFrdc7Ft1d4RJKyHU
W0LTjz/S+kwOymcm5OE1waB2xZr160jKJ9TMG8oaN9rnK0xygznlkwqIbrhcTz/Q
NKBA4V/jtp/2G/rzpOIW2jxX7xWP0zi5XRVI1GsJOHvcaf/NGd6nnn46Qq72tl5F
caZnuz93mgUPhzN6+VGr8k4ZcH7Qv5Y5r/26WZ+9bPEr7EjiHiCzug11YrXiXtzD
lU0TokgEiYOcrMjdaxwzImwQcIW8hVJOu0APczjbuEY59BjGTTNpGwdCETfJG+5y
kgfHRxSHy0FlBa/ErYVOnUK0an4Zw5e9JeIzENJDIzpXkmAELNSud1Gbn4lP/BeJ
qf5cotta0yTyIFWGBwuhBzVH4H6u4tOe8paCoMcJINE5aooMDGWH2SS98aNQ08ch
sMmfMlhlX1w3TUu4C5+JYp/Oj6DRez7TYJXh1UDGatqyUqizlOvCupLa/rCgu1Gq
PiC2VvAp1NnvuNH5qNTfGO0zDb0/s0qcOI9YkcjAPU+K94O3l7CNgVGjVhaGbKfz
1TyUKUsqh1huRmxWAEw3sj3aCXXh5GKTOUHh+wN3nWDxZhb2TNWlomHl7CvEBHtc
xerGVV9a360Cz8rCHNre0jnhnQgH+VILpsMzyNzMPy/hRYWpWuJOGrS2JLaTNx8R
q+K5J4ePJAk/kN+pFslKUzTiQ1y0OFPx63fs/t6OcQLF+pSKdB/o1Kqa2M1foBuc
64LdAdHSQZdLwv0lfgiX4Z4l/9hFPVZbvHnBA/oaHVRIb/5iUC1HAKAbjzcfrus+
0LBRlDgNZrKTcbbaRJ819w==
`protect END_PROTECTED
