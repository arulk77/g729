`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB2eF/bXHWoOAFU7yPBxSbelUuHwxe7N7gChWQztabIj
csXyJjS3gmsCaDP6WFlgP7CCue0yUYyZLc+5RB0IXs1GLSfC3m/MIPoLN1shlJFp
Qfc/XP9RvXwhYgk5L0/PNZf5UIZsep2AkskpxQ/4Kr8QfEF0iHqIQkfTl2PHeWga
GhQNoZHf8Memk22qQUSzjfd3xawCIfmljDZT9M1rFsspZul9vtbmQ3+2V8YWF+CE
MuJggWQ/wcjoiGzbuQc4SNZ3RizItq9TP90IFxEFBsvvMi/uQ1LG++UvqlGOSQZe
6h5Zpm/A/9szHj/wf0/IM8G/1oajBfW6vhs+/LjMoCPsKUKRAGCmvV32JWEpTdHl
DyRYCep94r64bYQrD7lN9LLxiuecMFSG6ErSyBe28L4xtfG7PBomy3WQDBZdVmob
5g4biVU/2uij2KIMdSQlQUI9/YwQgOQBJImTGuNBeBfoiZ/AZEMLegdMXVhmlUtW
La1bNHY10SRtdLgnuhS1GGus/HMZ5r6yrDeSjErfzwf/i31CtCdQNDdh/nWq+YW9
`protect END_PROTECTED
