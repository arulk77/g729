`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePkD7kDDUb+zgvpXw9UImaS7HgCyesb5PBvewkEI2Z8A
/1h97Y7vkNOQrBg6MTPykJqWqE9zj2K27JoCKKNIkIx/+3yr3aKz1TKhLVFWB9K7
d8RuLcgpkJxecqLxiks/TwMOmJLpMMVksyFcLAxQaCL6o5NpVLh8CYzyouqamue4
QFsUXREqsWLwmZZCkAi3REjCzjQSao6IiD72xnlOH5LV27mV/bFt2uv6YGN49Gm/
`protect END_PROTECTED
