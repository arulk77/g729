`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOs33vvQOx7/E/nXwIlQqILcyGrAODwiAUFwiFQihV+g
t1A4ejbBqb1/mRE0E9sS23P1gNr2AWoZ5RWuG1y3ardUW3ksqutWl9bAAYJeOsel
gMgaLbsT2rE2VnDOEMDGhnCgriebk+hZAEyTUvwIB/FDGeaQiBFUqEyoCFArs7m1
oXSZkQmIhefO8VNHBlCQqSD+Oksjo9VNjcOMy8FrqjbDHN7kl9ETPWh7G2WemnFD
Pk4PYikJEB2FjBt0mVKAj+D+obZGeV60WQiij/T36WrIlgsNonEBGLxeS4NLz/a6
1QmkYrxkjt6d49rAFNZp4w==
`protect END_PROTECTED
