`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLfGZ6mCQgyEofwaVxptMQ4nD4+GC3kwghzi/RmA/jUS
67USF0G+AciFopZOjzdJxkjqbU+eoFoUdrv0Wum1Xr7tA3Zyb8a98sOQc9fovGIu
RIiu3SKWrNL3PeJjwxAaToW13PjdCsA0j7DRYyEDGcA2mia4IsdKwpoPxx6ZIgop
hnnafl7OIC5T3YDAmK18WOxGW31d3xx5JXoi5xG+vM8wVDzK/2LoBM3kcd2XkLHZ
EOXNsu9IZZt25vAP+Y/XjQ68LWKAYoumYzyOcWmQRmeOVPutjwE+RLtKsDBgo5d0
83LEwoe1wf0wkSEDeR3wOOLp4MiW+IpzZw4bbaeW+VE8GUPQmiZBKzL7cn+8KFQn
HrQ9SlH1A8hw2RNlPZPcJfG+u2Gpp85APV6EIitk7uuuDLR1+dF/FJs0Df+Urq94
upQmYD+dEi/wBmiEX5TmW9EmpCY7YWzH7EJcvzA/e02I1l//UspaeBNUyaDb+Jw7
nD0dCCA63uYLIHE1OdbCtnv+uVDSoI7PxfuTujL1XCZFcBn/Gj4pUD0lG0CAxRZ4
7ehztbjmeBv8IXRJPyDYjxNTc/Gbc6Mytilf5KBIwLWsGA2cMNC5SSOVJtmIg5hL
vJNTYVCyefjW59mBiZcwPM2m407QAxjVusltioFA5ngiHCM1v5cP/TAHLM6fZh/2
C4hfhfzlQgCJx4Lcyp719fo3uFXszGDCdZd2LtNCWX/DwWLh+IaFvplU7LAsqTG4
VcyB9v2CBSgqW6n8js8ObbUWJq1Ak9s+zKX6Tzbr8UsU8bu2ttFTx3oDItomCZd8
3ZMDdAyN/cQPBFAoQ3LzDJgngGja1eK/Ct3ZYH22vKN/ylsDP7oQBOZLsJiegdgD
ZCS3Ro7TolQXzpbKgSgBD2Z9ogxdNWSUeKTeyS4aESvdbtsKeC5yGxiO6nFJHgdq
KzJakedajXB/oX+rD9fs7/RJLVGGfHgSppzE534MPvWzENtkgwx+hRT4NRWR5+b2
`protect END_PROTECTED
