`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pLPZfgJqiHUxNiDY8/RKHrFl+lKgfDY9q6Ok0FuiTOAC2txKR6rEM687xJNhnKH9
yw5/eU0iu+b/dbgHJ5bSAAHFgJNLiJd2NtLDrrG6aTruZLQrmGA+Dl7/If2gO/RS
qrBVpbfDdXfAVDKJ5TV5hfVVq7uV+/A6J/OH/IexqPxSHiQpMrUnbIEM9k8n+C9m
tImHrGJ80CtiQyJLUAv3ddaAGxNkLGW5c6o02SZauxfEcpTbHKWcAPQgHAgLpnQz
5VgHjFuD6xsM1HV/z+cdFjiiAd27sNXCx+YOm/QDVvQ/SqHtkPbuK5Mm5N2Nxa7y
ijTzFsr7IJIzjIoYo47FrqviQC7wA/ar7v1B8alODnjJOZb6Jcw4B0YvN3fKWtRV
NnZ0Wj+wpbO0gKHELlLSW+XmUGRjLaLv30ezQFsmG5HpzEifvR8jt892v62D2zrq
jtZ+WaZ0BnLHa4ZYqrElmbnr94IBwXmC3wTb6gDND7rUT8fBcQnYm3g9HnWfzaKz
N72WTZxSHQFcP2lVvAr9QTuxjZBYCrD+H8xnQiknN0s8CeCS5d4mhc3btwIcjxHK
OeLz3MgfhnQ/R73M4a/wV56QOGs9HDiqMM7hXRSATONN005UHhPdzTLnShU6gON2
UeKssWvGXlhnoeUj2Tuh3nezkWR4viUZrAgfxXAgyt6xHg/1Fy/ZeiR5QKVzWkDT
tDBWwSrd1PNgHRWQi98LJTSGi4KCyMvxiniDGoC+8wO4KjcKeJ+3d+2lnifr4dWS
kj33yCp6BtXdrJO8P3LVIHOAEkRWerEj/92XHSC0mCGqmcy/vf72HXbesB1fuMri
UWIlIX2lsjTSj3mAT5DdnA8wgBUfQwH/usSBPNvbcCQSpT6lapIts79uPzdpO8Gb
MGrpQKExU2784tW1PC2r5lWyYqaJfYwGZZlSwxo9nLUhGegxL+HfrbGUZ8VljVMZ
9pFFIgSBVG96oHAWZY2CA1h/bc0UU2TpSGYDTLYor/eBIFFGvA8EmpRkVq40Y6aK
zyFRGEC1ixcfnWDNghCcWaugNGbTdVraTUTTMPzZ6gdWt0bQhmV94W/rhr3WaFoj
yEuDNKSDsZDQe4Cx7gyro4Wv00PtLDt4pmo9GU1MCTvLMMKei6cQ1utzz/ihC0yR
gzhn60Eo0e6LuDoJmzmlEUvfT36U7rOFnqu+3EuenZDS9TT3FCeZbqUr74OMEwBE
oRnYqP3S5I3su/ZKs3UTlF2bcOdRZmqKqmqIdOkJaOmcRzSzer8CcZH3xM+C71/y
WFCsjlOBCEXDGhvFKvUftQGyMlV2L8TxkpxiP0Hm1TOVJ/3DrsqSTJE/0nYtO17S
O0u8vTYv3RYbUUSh6X92aex2Q13wMGsA9jNrGj32CzqpE581V8bICYnjgpXTDd8o
huvqwPe18Jz+toN+xS93cQqkvqNDaDp6h13WD7lmlubdShQeunBCAk1mN08xBRNJ
WtuXO9u4T6D0nPErlCU1BeThhZQbG3lDfK/fLdRWpCSpBlneEiQkhfRmUw9pssFP
sY6hNcAx/JsRGyGwotAPSEqaHlClUAhOkVSE5+jKvfgHAF6OpT4aMtUZRDimYaBK
Wcr9JlmYzKMgTl4KN6wLcETdxVWRV8jpmbsExFfV6lWQkxK3wLciTUE4DeLLucJ6
R5GekQo6B7O72HADW1HURvB61wyS11ofO+FksiJZ09j57gy229ktqPWNyGstQsC5
FTyUuL66vbUERAolxFtlSnksoc5c8nIqN5ilVPQ20NZjHmXXQcmrGwlm6SfsKfws
3wmcVwozJ24oytAxyK8sHjV4JHlKA5wd7Ncs7xHoak6JeZU6kP3uny1L3u4hWmLa
9QUW5UNAErg+1A/cLzyXK95l6PPlw1JaNLA4cG82nEPo8GiNnabVNUgs1P5bf84w
IEejlVYlsrjUZhtwtEsuvQ20yAXJgRIWtXMSB4lnqAv568YcpM2ePPiLbQknKBUM
UinP1lCcvx3KfAJX16Ug7FlwulSNh7o3weiadLemzRqV4oyaHyT1BX+OvQ8e7b97
FmKgshFZaCXEp0o5XLMKzd7Eu5wRv45+OFuntoqmixtX3P7brJ0lWCHNZl9a2p3X
dGAXSMtWJQKvh6Qhsq71UG7DqagAQlXGrervffbwM9qQzDIM6kNZ9vu5p67Vs25i
j9IPG3gKOuoWskqpVe4eLNw0t4n+ZaX4qCHGDhaf2JvycYiH9Mib2fcKs0Arrlrd
`protect END_PROTECTED
