`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIl4+D8Ot1728oqguMLxWCt2ahRkDdSSv2wWGSxDq12U
gcDDpnvrQ+Gec237lYN1QotPKnU8x9P+KCB9+rSSYidC4lEx2VBQF/Ajp82l6Tmm
ExLjdsmOe/+4ai80O3lFM7KNnvAfyld0nGmf+R5m8hyXLcvuKRANwlztWhlzHHVV
Mm5cMvVXGyRh9B1bTVYmaCUH27k2g6ImugPe0qkW5RdHFCrBHPPlwR2kMuM9uHVO
Ek/NQrTThPj69TEEw0yqXuO3ZyLISm0I913mY4dtLbhbc6l5CcCCyrSdou74utuA
gcxrpIxr/b+lnD1wr4dJDO8mO3zQ8tZEXz7T47pqIiz7d5t5HbNS/c2Nf7DXmhn5
6arJjx3h51ccAzLz+j5m/SJlpjBkv+GSsUHPMPzHVZylfbFyvYBVDQ8Ugei+AaSV
gbtlZBMfUnAnxS/QENdIpd3Xmy6vMy3U/Q7KWK2ERgpls0snt46sTZjYHOdP4+y2
34s8q+APWmV/PWQJwQMd3iOkp/Q6Zp7XlfjbLgp3fTKXBCLbRtxMRdDqzSM61lVn
`protect END_PROTECTED
