`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
d67mQtZ1bv8AXNNz+L6obhXc3GO9RQT/cLNLulLm9QoGZX1JKzYZsg00BDUTQIAD
Cq87d9lMl51XS+PpAClJuAFU2dxDTg+81DjpibCuKiY//cf9HL/2UDUuZ7jW/1Yw
/WjXDCshAoMv7c7mteDz1Xb2o6sulKrjjsmogObY5bjZtWP27WbXVSjzGYkVTrRX
`protect END_PROTECTED
