`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLG8a6DmMHJr9nL+dwBew7OaJpk9MGEDc2lgpLCHBVQT
vbbGHLtB7vUrjebtIimSDyaKU+RuiSwCbqZvZbOxKJX0Gr9NtFo7z1JG6KBmNFIV
Qvnh+26aoh4Hcypw7jGHGOT17i1Rig2rb64M0N1ZOO89bR5ODsmXyMOjVYq468fN
9SlbShs3TCrcCDKeVaG67PHEoswnHq0hOmBTatpuqHtp3XJkjCWOYWuH4diiwn78
`protect END_PROTECTED
