`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBP8GPvnU5azx5h0byDhD81IRBeEgOoRPnSu8X7Ss0pm
VAmcWrmDDoxcl65TdEkr61nwy0pQNemjmclDBKJM6Ewzi8i1efsZBSzpPcweqe/+
6jzUvOWDt3Lnf+wudm5F0a8wS/oun3FAFai5xa2fkTwnQxcs/kCmv9usCq/TO80X
CstFe8gDDYgip2TgErBLgAk374QwvUPmHOFbOwtkXNjmyT/1rPUAi7v7oMJxQoqJ
hE3Sm3IqBaRpsKF/HZxryVtEQjfSano4Ottpk3Ypd0O/OpkCfnylEMiB/y9Sy1cP
jv4KSEvuLHyp+sDeZBCizWtE/YOUPc5Dynr9zdobPYS527PSWi8Yc6WSQ7dqUyjU
OKP3+ncHadcERE2cDLOXDfO5jJvlgu12zpCw0IW2EZ+xEt94942r55i/Mj1lRAz0
ZPorv1ZOc8XBQfue+nFOPzgmkOsxuHy3mFCqbLf1is8=
`protect END_PROTECTED
