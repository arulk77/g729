`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
g5l5AyvBAUjVYnb+CwjhLSFwaNiVidXifUrtg4nRJVfHTUu//yW6pHaV9UfJodEe
BPP5z5kENLKJjLO4rsjAf4cmAc2sEyZk+lt1D3hTMR2qYrQxb4O5aPVACw3HNUAS
0R80UGngrA04vXcuqxl+aoiFKsG7EcS/lV7vUTPi7ZDJNt45Rn6FWaOGz2U9rMkE
b2bt0XNbUqlORR7LXBiQsprYF8aMc7a+JFDmWCIBiRbuyRTWI8lCKsFM+xQsYtP6
l4DTN4tVXFNmkM1S2KsPGB2Yr/eKMBTe1DHMl1jz2+bh5YkgRqz1NW2O0iqW8SAt
IdZUc8PrJkHHnl83RPBkmmRpdme4er6l242/VbLCgAk=
`protect END_PROTECTED
