`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDGSIKQ9JFPBuSh/jGTyUwwAiGZkixem6+K8qJesZ3x8
hOBbBmGsey7sKAiHY2fc9W5p0ca7Pv0Qc99PxwRt7UCM/nObhpPzUr1v9JN0Pto4
MdqeHEWaoy6emaypS7TnA+Ih9q9Woz4v3EbxnvcdAhkpKr3hqr65qsrFms9rraDC
dBu1p19KPEZNHxyru8ggw9EGIC5ApNgm7UTjc1wxGxrMWt3cpnjg/ORiHPTWg62r
fKsnjivPO8WPTdLDsW2t5dUBy9ZLtDnwmjE2hlwWBJzTC8Y1zghv3A9U7mOzxtIN
dgfzjOeHD80HUKN9sWdedJY5VQKxogfXlimdUggBevvEIgUQj0AG9L11fA6xVDG0
hAVrYQJP3zhue1v6flxoQWlt/wIV77KsHEUqVNJdaJYspsz30rAIs9FSX1uzx/f2
7QGFA6Cdh3HASFTblCg1DCJzHLi3vVxyTH04LPu3rFc=
`protect END_PROTECTED
