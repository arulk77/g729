`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49W7hcxCwqH+y2LImyJYmsfQmhUm1kB68NDDRtU8aB29
rbN4dZJlqq1wHCQWXoZp4I/VUX5BJSX8RDZ7rey9xfLRgSunqumG/DZo5fFqt0G3
QrmTMQZGABa4bJp+Mz23BSsDf+nhW2Si5dicrJpXOOZP4s2ywieHVF1kfrQsDWct
I+0BhyErhsFYm88vS7m+iIo+i5Iej4qprwjUODF4RLyefXZEOr2M2+rRvXuomKQa
xG4Xz5cijIM6Nu4JUBC2rhyPmjkzn6uKcZOV8VaUb3vKUV6nCKFdMo7fh7de6Xrn
jVzUPqQB9lc1jcLnTZdrsg==
`protect END_PROTECTED
