`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLilqBf/NVMabD8GSaceWRsYoO1FQyQWrY32U6X5viiC
90n0zUCIj0SspAAKxRltmyWrsVqqqwYN1l6eGNJxNwSDbHkd3ggGDzFsHJfGLsA6
AcJ27NgvF46TZY7S/JOoocEx/Cbq2XccLq9C9O84iuES6bbJb6ur37YbLgiYyj55
`protect END_PROTECTED
