`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jONFBO2xVOhASpI0W8TY2MABxaOLvx2QQH3FRPyY1LoQZ8AH7ricUJKSeC6Gtkot
9v9krKXDfls6PRnJeaf+M6eSLYHLcxNHO0627dWOV/x7QzlI+kvc/wYjj9lJc8mT
mzJKspGaSq9Hs283MVjs7U/eFzv22bwxhb9eu6LV5yIK4KE+dPIgp+oDuFAgPJQ0
Bt39dqWL8WnsmuKB5nXdJe/T7A2Y74dm5KCuuh1sCynvRou/VNbQQFrbEQ7Vmvdb
9T9fYRRNiScpfllaXkap2HYZPSDkn/hoSdY6lGgcCyCrUk8LEwE9w4K2UZ0oOxmM
CDv6Cg340Z5zrpwrYZGf8njoNBZiX/8+aUluh9fDAnQ=
`protect END_PROTECTED
