`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLk2Wz+lAsKvgava+ZTI/0F/XNHPIgnsLZRQLyj1up7o
uK/wafGQZXs/hnhINOA02Fgact63AOZRXq3rcNoXM/jNbRmSwPdJ/xyyalqZL4zX
sV8lxHtt2n2I6xNgNq1IUNsjADsx/eLVOxpgQW6owdMs+S2Ktup0kx6IGAh+2tHz
WLm4+wkXfVkNpI2hZSW7gl+b1ZOfE3HxMukIXQVFaDbGFR5wiweXa7avPdmHaePu
1QzC15C5YudNmxs1fZR4iknIS5KQqicCy6nbc2MQ3zatH7CO49Lyiu52T+a/nGdd
1eQs1Sx4BAmrawn2qRtbqMf1DGrLq6LwFTMGkMx1p9b7KTBM9A02sNQ0VBnrDl4C
Z0IIFPoC4saJX/CWICDUqspZhgc2p0nzEeQ2ec8Tyqs/XYIESYAcbJgTraUbSKWC
GpTY1XCDFDcXLFkUqkQPfwKZ24BoF6I1C2gdx7zI/U0yZdAmTEToFtdW1oPAwHLp
`protect END_PROTECTED
