`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcIDslL/rSBG7VPGW2Ssvflpg6NLJqNcS1l9nRie0NF0t
J/rUQCBv+SJ2IMEtLDB9yraPRvjDzW64qAAJ3sq1UZw4Px+Ljfc4D7hW36PMnYGV
pmTOusqmesQq7DJFPw9NOX5H+de7XP2mmwQSmnUFha9+Uwc1Z06CB4FwHLvl05Ca
qXOETGUFIO492d5TREnGEUFl/8t2yzfZ9S04X7OGPu/slqolsGx1QYDHakeTuMwh
OjzqH3OKsRT2QYzMfrboE7mRS8+NX4y5cCgCJcANUDew8VbI9Ou+qP2JFh+8KOAu
JsU5EjJIA3LdjQ2KQ56/dYImLpdNgeBZzxoO3s3FgFh+IWU6J28SN7qGdfoejUce
`protect END_PROTECTED
