`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI7tN3ZnuA9BMewVvv+kbiYhsY0kkt4Ny2E+JVSDJd84
ozP+/q9roU8wed271qN5/dppe92gM98fkmW+FO+JOvy6BDn+1TCvGuZIW7PceWcz
+2sW0rwbk/FTluVEH0tvCxxhRuYoH6POoBMOZM+l97DMLqSBqGG7lvgd/HvOTxf5
I5CdG7Sd8ec3vJhGdI+0YVCkG4Inz9Nt3mlPMHtQnBpsyGYRr+hD0Mn710AJghOK
`protect END_PROTECTED
