`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGDglPWR3rC7RiHQAaX1kQGF4clfQefnRuuLbJo4MHov
AjGyfO1Dbsj5K1enDvdad2xlAuH0DUzbjqP1JSmYZSLIaL06Y2lMr6YY1mNMLN0r
bIL4e8y33B+ANLoeJwoTyw4Ce9RDRhuy70X9eARTX6q/kNN/9gzba/gYGZizlF9d
xSN2d5NXfzc3bFV8hJSNly/bzEBLXi803RI7JKtXf4FrEyUMIJxawKklBDh2TBn1
/cy0eXHvnZecWIUs070BHsv81pd9cXk7IsX+3gfGPOjmpnpO1BIwsUjkby90xX82
zYWr9Wndt+L2qwjCxrcx551xHsECeVPCH6uZrY0XxE12mloMgM9Btd/8ttxbW91b
o5Z4CFv8O00WHrT+3pQ+HbI1vSe2FdQc7OdNcgOAtwz6r3eWrgmrN0EQdz59ezC3
L+SpPRm6jjX0hqFZrxSbR1GCIcn7/asXFqjDHAQ5LGZ10m+zWhBl6wJ8hdeyvhTP
NUgeOvI9NjMVUfjEL2rYFOuyrQ4DAeYmuoBj3UO08mAK2e078bHa+q4RH0sl/CRe
m/0BuOxGcQzRnNEcexxhNwWM+aFGyhb0BDGnb5rRwtXdqUjwxzc8Y1GlSOWHaDU1
OeFXXLmrwzooX7fc8PTkWbKxHz38yOraLAo1XYo0Dor9a8HTbDVfJtCODQHHcyW/
`protect END_PROTECTED
