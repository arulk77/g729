`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wVVJ8hPgx3Xyq6kosqdkcCmIhPu1A7EYR05RSgETfZP
NA4W/ilMTe8A8isFQ7uDsfchWDrNx4foiUFn4jsJw9LhMZLmiuDB2LdId9UWbSuf
x2cj+61xTFHVUq7MM2S0huOzB5W/3vP1OFftTSiD4iaajmuXJr1kb6VtwjqitrMJ
sAXMHK6u+F+k94KXZpbMuxzvKILJAT4GVvbwFqySGkFXPzErwnVb/cUBsFUiW8Js
fO0F8CUWWdVrGp1zMbQet9ie8smcNS2O3rCdg5lDiXM=
`protect END_PROTECTED
