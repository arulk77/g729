`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UY+0toA0b0qRqD/tz4dWVkeYoqeTMfIpjvaLGSPzoLetICW2GMVkCgJLZSKKa7Bx
WytcQzIecjeC4KAx87FOVusRBpwPTUzOzRzq2wlr49jn2tR8rAyr24lviv8ZLMeK
/Z2I+DMF7qaPmix76Ti558Y45q5V9d+Exc+lXdBi26BTXQfGw10Vz99vwcSNtdxA
IDqh1YH/4q4vqi7qF1KTocRTG2d3hz6RYQXf8HSjFlk5zREz/5hkQ4A82fLv20mh
`protect END_PROTECTED
