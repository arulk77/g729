`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
B5yip8e3mmFnxVC4uLPsDf0WxYj5ZUyinMcGln6I+wHbbIiTaz60BDQrkaxMwWlD
Wj5A4FRe4MFFDiaVDrEdCoM+HY0xoETOG0mifXh7dyxCJ8BdK/ZNtGxsvWoOV9bN
nO4BNNnrOOg8ao7Oh3lRUdx6+QiMVew1yEG+RfqR92m2Xo6HCBj2vR7NuS8nT3JA
akzHMmod5AlhQjdvYcKP9ipBu9oTwt+jxKbRwY8/Gy1clWwTzgBny0ZnTwVm5i+s
vFcGV3OmY6uMqDv9M3rzaon/PbsoqKJdqOdjKgZbfFPqAX0HI/5mTekpkFta5pGY
sLwNDATUIkId4UkAv6hsH4+8Sxg4DPSiJg5ZnDQBzw7weCkE7YYIe+sXO7RlNQh0
UO4yTCdeDLanQeIviuuGiUOSDQxQL2GsjvPEUN4xHBU=
`protect END_PROTECTED
