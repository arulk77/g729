`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YIIZzIfVDdX2qc8vlTUQRMDJOuuWYrUCWPft2EiTCd0y751++aMsJet9vkwZv/Sh
Y4PiXD4UlBOBOyazdk+2CPFj2bD2wi43r/vje5vVAuJ+C2wS11cBaZU3/01x9o0k
bnHzGQBu06oOZp07NAi1ojCj/cvYqgtNUAbNBe5g8aJKv4hyOQCQYt89qlH2dISP
JOW718Wi7IBU4RPcT8I5sTUVl3zqR1DEjbRd8muM7JvPjj+uFygmnC0mSNP+Vtsn
IgbEvRZixZKZuM2yJT19lYb0LpEy/pi9TBMGd7Y2nqUM8iUgaoq1SwrVueVnHILm
1Y6AssgSWlp60njW0OXvRuqtc+T6JrvDOyNmYoR8184tnFVIPyRxiavNi1dcSANP
TyhXAuXaevA+EknvFnyYTGe6ycCsJjpVAktX6Al1IHXiizf1xquV39lF2PKagunn
VDUAJEHrj2iczVpVXlJ83Cg5K3uBxAM5o7MMDZRY84I7eo0/AfcWjEreioDw5He6
No8m9xJGiDUFRXMHzZ3N85oRsXqoFrzPPXMg+zAEjbSeH8cQEdXDR4c13dsY3taV
l5Q4dmF2yM3FG1iDGNXmHCEt++ZEmh8kQxPwP+OFTvedZstd/vIQkjFe04zqArVA
TtSpQ0+XpLY+C7eh0f1/Ww==
`protect END_PROTECTED
