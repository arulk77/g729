`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJK3Lttn3DGcJBQhQ+2q+2NPDkvvqDjk6kSSLCeI0VRg
mz3IrXJIFWmvj/DeJvWtp+b0p1jFaBihSTKcV3+/OrIT/ScS64EPCURhPNGiWq39
h9jAWIv0QhIF+G5TcoqkARVg7Nlcw/WKnKNmqzfzj2VgiZDKHBh31bP/+aFQXSkd
ruReiEuarwez3Q9X/lD+UQ==
`protect END_PROTECTED
