`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNye41YMUb+729HmTO4oXa0WYMDMKK6Uo8xmDECMkVM1
mmFwmw8qPHEaPR1OEYOBiN86iq6C02TWEcVZciGVrTyOWSqkqLk/xWNykbFaP88i
bVb4PoqUoDneCj+DJ+PkjF5JXsq2ev9ZmYUdLVO7tamNNArTAVaKwn5boRy7mn6K
WASG+oxYPCGMQmF6u2uR6HOSCFTcOMIg56H5LlW5/KOaNObs6ytWNQS4b38pJ5DE
yAPnPnta4T9U0AKAE5gZT1ie3NTOrPQjWZGf9n2GjXbjhSZXEyyf2rygVh8L8Lpq
D159IT6dkPwAWFh5SzS3xyPcxfEwMk/s/w86g//Eljxlg9D5HXmSUMMPEShlg5Az
szsPibAQ2xWnb3Li5OoTu+vBL1kaLk6P1f/QwykZSFxRS5yHkGljA7b7Jv2L1VOR
1aysoZgYYm0z3L507BaJrfdDJzqHF3NqRzQzyyXTfJGbHNXTq0Z2mtF3v4nlntWU
aC/t0AGSzvpGUqIRs2PS8Ii5ha3Q+5/u+e+zlx3yuaF/6BD7hC8WsE1t7+Wfxk4W
bPYI8r/fYUJNzGaWLAgeaH0DFfW8xsUNQHOv7RrRsmc6E3vOIb/B1t8yykuV8+z1
5tTYAXT+2w+XAW7K5FICb3di32r8U2ghICdCRP6J0hNKeDWNBxbXjDf1/IxBNCZ+
`protect END_PROTECTED
