`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePAK+VsgS8Z8brujfxrAha5n/qQXFKUpZjZ+oqLOlS1P
xunJFSndLg8gTK+btDEOQkHnSpsC/K/z2OBZWs3lSb0ewYGs+/oeY4Sh3QVHR3K/
5JIgeHXJ+lL2pRd+yHJ8zVxvhuOOjGeGKUB8+VQRuaqtmyNLSSUkE4vCDZXLoP9w
87KGKhuqPOe8AxwGCNwmDWqjjqG16nHdfND+sJPj1gwpmvI64Rzav75aIqOX8SI8
QCN0ELBZfNjSPRIq7SqJr2LkPtVw6XBAvYvkQpG+OWwv6+3ei0DAuLC0G0f3sHI/
QA3HHdfjb9pXC0lGkpYvZK0sH9FpF8KwlbzhcdkrDC385k4mQdoF5fliKMuGBPWl
Kqa5/JtFizEssxUkriX1RhzZlvFxWTnb7DTjPXm00z42SeX01VbruMqDnkeR2Mqr
mhPpqPeLcSFWGOQtvr1dWtsx9jbMpuwzbqWTG4pi4WF4hPltuwy+QQ0FtitYhH3v
8TI2JZJ+FabqgvruOVUWwmcYxZYvVrK33LwvYL7loQQiHveWW/oaMrdcjlJDaAWs
8luF2UHIHt8LTc0wxz1jmC370xbq5Ovd5K2C8pkNTCTJaS0NmjoMXN1tGeQb+PYu
vw648hy3AsMpWJqyV567NtHwPaWLzNBxZlbVu9+YMpFOj6a7RoMRsB3shtF0MXfi
m5MR7MbqdiMVUAIzgUXHY2yT5WK9ag0A5TpIlki6CwVFM7nfHQKYtxzeB7DfJ4Vs
eF79/BObRsYJ+6sfKsfLZXU2pktPhC1nMWuRWxcdve8=
`protect END_PROTECTED
