`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKeyi4zv4hJTQm++Xm07bIe7UlxcuF9o8dbNcG8sks6c
BRu9MCQK0pCgyTVoEZabLfrtfsj32kwhZVzj7TGB4RNxLhdNWd/YwsVOr3feolwV
8Fn+4zrL/WuCTl+0D0V08okXeHb1tgwt0DVlECLZm5zS2QsPeSjVGt6grCOJKgX7
EwUbuU6l/1NgRIjuOm311NI7L8O2SU3GeHQpIajXvbhUXk54RMs4qaITnARk79UV
+oWR+4QtCVeKDFw3x2UBcw==
`protect END_PROTECTED
