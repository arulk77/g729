`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJsy9mjSiMvDYJRD6BqxDU78Cq9ri9w1NOhg4fJUmUeb
mMa32t/P+I4jpPpEAmn9tjk1p8f2KLyFR38h24wbZMFVedjgzrgEFlPRElUtCkoK
cSSJBb8qLSS2BC51xbm8WBHSs06AQC0KRYKS7oJ0cJzhgz+TfQBv/cZn7bnCjR2Y
birJoGyz+ArHLSExlqBv+X14nYUHAgg8Qd0a7HIYhDHhAwAPgxF0u1DhWtac9p4Z
U4E/KjyFiJMqzpz28f2JN28Tnjlt2rSA17Ue2sZSsbH+Y0yC3daHT25vtyRxXKfN
OQUUw5tyYK/DxYOQyym6LfM70qAK3XLRKpDup7Bl7xSHuVud6NNg8CLjayQfCEoS
fO1Ptpe63d5PGySS0/z+7Sk9LM2hU6TEHYuIIFWlSIsWd86fBcuX7bE9/Pxc4Uz7
LnRAYn/uzXc/g7hGtv2vwwaKcVEwK9qML7Sk6S8RR6gWEn0QXeRHVZTi3+b1c5+a
E6qDWynh9cEOWQXhZ3Pr0gCjX2tdOIKp/oDYxpixG82frNnJkihfauCMhj7jgKho
kgd4AmQnSkaoUWVPpEZ+57UkeoaNTvSv4m0Ru02a53J6RfXzSPECboPr+ip2pHTw
`protect END_PROTECTED
