`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL56XbzHEPPHfH4n/5NGxIt1bj66Lo3MjFS+6jGoKX1E
+RtRTg9ds3fMneKlcZuwHdB0PSI/hNY2dZP5QGJKmOutMQEjK084aRUlCbITa88i
DMRJF2ql33PZQXUyzbkHf6OWF1TV2EybJqEsD6rxLFTNbtj4vXfId8xYQYtbkQ8Y
TOcxHcGNLHeJdSNVKk8eLVKHk73HnpRYCDJIG0ls4tGvrGgSQf9pFQkxTi3chV3V
VyX2aCGfUCpEieLNvN0cCsz0+dzuzxGpezH7lpnXg3ZLgeB1O84xRrvjvlKJD01K
tYGLLFGp0ZOqp32doIjR8BeRpJzb9DQp0cn2NJ9b5BTDG4nuwLkDn50mF++taqEp
zxyPMsqpCQQiH547+vuBsVFmdxiyBpZ/ieYzC5WazGmPdesxjn+xGXjfqwD1ajZd
qxwHYeF/07LRwJ4YerlW7sF4aQG5QZSEyWf1MmEwnGK9/At2tbxkrK1MStKcL5Ic
MlFEumH8wwmBEeD8H9yYwlre0T4ycr2gZo3YAzh8vOMO73D4NhFMySgjwiJlSjIe
`protect END_PROTECTED
