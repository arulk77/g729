`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu427E1s8tTsDIy2yRUMgd8IIqQkswmSNUcxcLYXLQjGzb
ktl+TfUlGORsH/Q/Q+4KvJviawQyDlqj7PRGpaUVccH9ZmzAeAG1JWSNZF/vIeGm
GHDlS3Muhi02XP7nDzLpkAXGJyM+BRvkV3WyOv/Fe/zusE5CTC57mBXJGWiwTKTw
O3f2kb+X2IdwLa2f2ESJoCkHT58YfOjP10vBEIrbWzRb3pw7SKgWmYQpXr3X+WP6
ZFOLceZLZQ1dXbpMBqhMo2T5OpazwgrMQvttkbXiosIvwXiujvXb5ZHTgax0xvG8
jbek2GUlV1EluoBz4qxBC1wFdWQj8tbMKKF4uoXfscgRr2B+ekyuQYspwnBMezYd
IeBxFt+1byBTXcM8QOIyeg==
`protect END_PROTECTED
