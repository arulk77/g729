`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45CvrWV8SdAO0UT+x4MTZUprB/BITcPj2JHA2i0QqfBM
hzMTk4sE8yeWXnCWEGlVJfwzWtOPyFY2NcazhtcW1SVUJ19mjM7C9Ke5t9HoFQqH
SDS5Ib0qwBGsNk09TYOBJ/zkAKGIgCB0WtP7Lgq3J4yhSqzJrAw7Eyo4NXYsycgK
cEBw33cOQSsE78qQn6P0QyJKy4S08Z0PYIPGrGLDDDc=
`protect END_PROTECTED
