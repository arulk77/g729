`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB0WO+yJ1vy1fVtpSL/1+uwnh/Wxb7wAo0Tor6mhCnxG
xyBf/ubUurun3XMM8vZP3nl179cSD2LKKVGjxdYmLUznJT2QUXdVCUda+71uuOCf
tDmy0YUALjjhiFuD/toks9hbi3EtQF/f5OmmKQw5Y1GbmJtLf3snLRHToBOrf07F
BBAhtTUE+cjAbvkCBx8Kjg==
`protect END_PROTECTED
