`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
d3BnsacJk6yESnBx3KKM6fK/z3PESpELVvTZhaWVYGNnyX7j2Mis647GzIBLxrcs
zhpN/zoJijXOt2mtKR3ZJe7InjRy4s+tTqdN5dVWE/7qmAuQhCUbAaqgSF4pL4tr
df5mIfc7zHHLbnRJTIj30VJXq3o+xBISsoqbU2URltYL9+fHAJPIJ3DB7yPmsM6X
RyC74cKxUiKnjSU9UrQuCHASIxjVhKi6t2SU/41HhWABPPPUIYa/2TjgLMOkq/3x
4u0md0g/EfGt0RpnWgcwgpsva2xw08Cs6dCiARQASvR0BJ57fXjGGzzFrmDhD8RQ
`protect END_PROTECTED
