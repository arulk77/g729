`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jaIvzHf+RrcRdQAZqG8EJSJhuFs/YKpgwUsDeHq7HCOpBVSMd5YY9SvqvLaL/TDI
O1tUSoYgdquPZYRPytzxY8Rut32nKzW15uI7CphzT5suQtfF6scfhir3iFpIXIXh
AyrtpA3FJn8Q10UwlqU2/EN3HvyU6g/B5mdTmKh2rtV76tO9B+xP8SpvUG5sL8YO
iw1Q7h+61+jPVrZ1Z6LLCeOePtgfGXxmGgCb3cc3PQkYPoBA+vC10pBO/i17KlLT
UkzfnI/EnjPTNhQG13L67uugy1ornrhkiDa2UP//zoKVTtHqyJ5IAxRs2BCV1Lpi
0j61wHh7JhxI5J5xmDqyVzC7rIwRZynwZZyJ5qHFJRaYIEGrPfkXDwEvBJ7M2EXV
+FMY8d2kI8LpgZ8XjswPw+YVkD8jGo5uHV1zYKMpkUaEjp9GAd3Tela1x+C0w3p4
W3YF5tLJB7BFyNYJBzrwIIUEzcLt6DSZYvFoVpsgDtZUvn1GudXskdGi7PYgeFRN
4GiV/XdJk6lH3Rika8hxNDN4cGvBcUrBMI4qWRXsuP9A865j7UPAzOR30da++oay
Cv/s3+6ljaN42KRltEDuj2GlsOmwgC0GaX1A2t3M+51sOAMRa+OLIfxVcnsymEeh
Ut4kTAiSSkLFrRo2n0MWCtzNCZhCF8SMoXaIc+HCgO9BtA3J/7cXwhr54VXiuJim
U8CtTSGsuBtn0yEX5MGkckFE0n0JX1+SwWIxQD8LZvToKh0rzKY98ZGuq7hLvB/v
ieoS/ao/4dZoJHcv7/uqVxBUuU7UAPu0BXYYqQGdrpFzDtFV0j05/fOREKR6HEXa
kHOk3WK1GzmDzULfsQmNV6XS+REt+jhmWU0kNdGLK5d6PrKZ71qH1dLaPgyd6k8g
IPzOYT5Xey1puo35Uegj+bw9f9OTZSDaRHWJTSQ2FcGinvd3aHWMmE2R2G7bkEll
U/glz4DYH6Kx0fwPQXNGDcVo7f8+owGPa7GjTYxhENfOn2n8mkpjiKaH+/e0EYsl
Q73YBDsn9LdQXY6NJwFsb+EluAwQunn8dNsU2iqWt7LluqpKJ/NWzmYngOhPnOvX
f1T677darZLsVarPBcIp0wKdwR4S1kdfcMY5ponSH675J3gXRZ24ab5LdVaKcZaa
s0BfGGPtC6iWmsPzDbHLbCX/Y4VEKDH/bkZbnkpDgxNUX8e4b6Tobdnvtsb61Byn
ZfMZx4J0dXba3jOIEZmUiPBS6iE01uIkhbD2Bhrpn137l5aVhvL9+oCee2qI9seH
g8i+AYBh0kAyQIBfFZhduTZ8bZWfLHTBeGcLcjM3QGUI9KiB15iUDlXhenUE9srQ
sHi6obN9Aq28AuCxaw0TqA03O0kbX8bJL6h9fmFM4cFmObN3ufaAJHgw6JAkEkoW
tA2VZ7aJFVKsZiF/Mr7qu4fPWhHcpHU7MVw0fuTBl52dxWNj+3hdTeZtDCzKzw3R
zzYEdWUCU4v8bNB0Za5taV/c82JeKKavh3p8rV2KgbrJ/+Gc+hoiFVABG3mgJhTu
Nvek+RiR3/1WJE7zPFjY7iJQ79FZQanOfUYYFQohZjPKtULioYZgXOvHRhb0q9Lk
F5Y331RqXfMVqd33dXkoXcY9T1w6XuwkGBB2C/Bem+26l6Gke1iETLjJi9dMhYfU
WYGh30//gIPy/AOgDucYcfTKLFwny6ZarqUmInokVdItHBnKeTJIw6FgEtcaOJXc
kT1O0oR8Q8MxAUjETDyepaypm3aJ+cj841E9L4os1H549WiBo8MZh/O8NbY3L6P2
vvlyFyRTkFcewz32NXtX4HVk9uZ0wymU/xGbG7P3C5Aq+J9w4oy88x23gUiZTs29
XYuLeVIP19JWmi4L0Ikj8AQng6GmQv5SZf12uFYhfx+HRbE70bGrWXsARN6zlsI6
ZmPHO11+B2IqT/6UzdlYWmJYxgaMjEBZXuh9tb4guMeuQtTv8Xhr2z5unTQI9rwR
RZ4H+OWThTh79iBNXk5IdpV2+dB/v5lqtEa9/+94mKTl789tCN9Q4NND4f2EA80f
OH13hpW5cOBHQectI5bpV0E0aJSb4MirHGi4T6IJE9J4wDCxb7tksBb1godNUOoK
Ob9J0ji9+F1NKYmRg0dGn9PnFujGd1+3876WHWRf3DQzNq+EK0VXAUuGyyZuh9ii
I1v7Y7Tv+d0HAW20TZOVyb8ffL3F614TmdoWzrdO86AjD1bw+QPAI9vBcB0gvg0V
dedJbjHeInOJ2dLcdeCSnONgvm5vlBgLeGpXlQEDGfygDJz5XMHRrZDsLbElHq/x
GFUOHv01UQfZuWSVBojtH/hreZsBKNONgH+scNVa4Tx3e/bpN0Exmfng996qNb3F
VRErIr8eWTNXWHDvt30xMoFN90LqM3qo96gA/fSqMSVaFCumAdMPOU+RScHXJ/gk
+UP2FbC6Jgf9zwT0tOOZVTXZbhze54zS33yqUu41Q3s8wPCiqevtheSgf2vzljA6
X6caS/ACsmPwsfB/QWlMMVgTGsSpchNUNc7XWAskE2/vGymAakdWFEdAcNqCV0oW
wLhlADJwRFAX5NeteFj4jpnP3l92D8dQIUrydKV+glTBrf3Gq7asDYSQlzP72Y6w
QNIaLq8iF1lROUvXG14HscBAYXWNUGVOkabk5FPd+7bEXQOlmfUak2l7AoJilPv4
RU09fySMQL45CtAc7/MNpMI0UIf0B7XnkqDU7O1bGbXKXjWI8+AFuhL56np9y1rV
9Tfi6qizgXyG1WL0F91VibRO8YsTlJG90Kj9xOjMHG/HOJocxfyZKKy/Up/DwH4h
JinwI0g2iIurBcGdMn29oGYtJBX93ufNt7dLq0OLdC/aRLZCq3m/oANqd/xbnANs
0yAqlxoMg8PRm77xVbcsMSIZxSvWljY9lFr3H8EWM3vfsa9ktJ5lWg9VNzdCj6l/
fFtkvdjF4VG0mW20n0u4yqAWU5O6ANpwqyTTB/DYPVJicrWgdorbBVfQxge/vOXG
hH9HkYdeLwayv41j6K8OYqLBOS+JrUVlQKJttp0OLUA6R3YMDMtc+k/8CbqlJfwS
JGp3ZyAtl/a1pA9I048Q7MSIyQpZ85HLQciCSKGRP91VKNlja/W39Tbd7KXyOmMe
GvuBAtKwuyP/1dEJMFu45bm+6DKCZq4G9z8TzNikHFFwv29g3tX107v3y7Ao78AZ
z5xfbJ65nKiUhDGB7hcDaxMlcKT+JDMsx/XmTovp8WpFRCp0tfDSfr3PKP+ZETpE
SF7ZsyXysFHWMNPoJMXQeCFBlfeLvAdyZenuZHXpmaX6I/DVlw4p8WMn+fzOTlPq
Ay7VUQN55w8EaEk9ndzbZG8sPQg9VFdA9xCFZBc4VX2aiDdJuY3o9PhwYagrvRh8
CFLJM+qzN+PPghcL6Aix8A==
`protect END_PROTECTED
