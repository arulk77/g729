`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM9oTLNh/ul8XS0WuoCF+EWV8DxIw3s15qN+sQclu3iw
gzTcODjCNujSRlZW2eOkMninYOqw6oiPpJVF2NcIEzK+0icXeAt994H4tX8irfFh
2vBEHdNQBW8wMjqRXsiK34AzbXKkPBnZZHw4Af2wvK1B7yX2ZcPztPmPp1fXl95S
qXCfSNHAwK+uO6MSwo4oOvdVRhfzOndSnb4Gp6mC9/LlXV364TcH+tb6MeZumV73
1rnkprsK+EhQv8PrStseKqwLG2q+Fc5W91mIKFpoktKfgNQdcWgKH4dr/QOEnq9O
FfatO4mCiJHS6pLg3m99qpqTQGsJbYSERotZM9N1EN1MHH2uEKU1Q1uLBW9pNvc6
N/pJ+0GJCJcmcslE2D5aTnKr/hWa2C4f4Mb02s0nV8V2yFuU1RrY7cteEHQj7/68
/k8dZWv9IXhYGdBCIgXqvOEQsC4MECJAW9h9nSzhEuUS/zSPdpvE3zwT9AQ66Qve
LwYUeah8XUBE6LTGdFfWeQ6zZI5sEs+f6XecvY3E68HQGwjYWXypzDgSVLdUCNob
KXisH332DAnHbfAki91MbME60/VIE/vDyjbMrSreUUI=
`protect END_PROTECTED
