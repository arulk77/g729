`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ssXPOxqXYHkc/r9612hiHI/O2RlCIAVFHfKCaOwqxlekqsvICEQDSolHNaZW7ETH
uwcnCSoNTNISPV6Q7SoH9xZsNi5I1oAoTn2QtzG9BhOpVE2YUl49W9JEvMCtzG/h
kI7GATIVbMQrjlbX7DJoCAXRq+z0dvV69ucHNNoZjqedfeqDxMvIoNsYD/knnn7f
dyIXDAFSCJbpGwlxI0stoy3mYyR1di74Mn6+M2hz8VwD5zDA+ktVE1RNtnCntlJx
6EwdK9D0lDvyjN+7gcVF8gzI5F0Tcieh2XTEAQKT/So=
`protect END_PROTECTED
