`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Sd0j2PfB9aZyx8vOrP2YmtTvDJnL4tilCGwYOAWVPGs/
3C3a67XjHCp1Rrwh5AWpGy1yY5zzO6j/JEUymRe1AvpuQ+M0elwtXfvvWRz1sJNB
lQu4P2S9iKHRwiKNK9gbA3oEtFf9n6mg9SRv7r+stlkDSdOewMFnlJkn2ZbPsXGx
F+XdM3VVcAW8dgpvpNu0JX5HDt0gaS8fPm4QWU/tJtAOU32ng1jEUoqyHjtL0F6+
vAdUcttHaUTYqBDxA4INmyWJqz5PVXTJBiGub3JD61PJAyHe1hXXrlNmbkOn2v/Y
JKNNfoSCQKIGhznicWxmmp18SRsIimZvedH8BUwyG9qf2ZA76TSt53X5ryQ5e8jx
ZbAMvXykHzp2P6RJLab8V/0HX7wduCErjmh0wr1fM8SXJPghLaZfCpOWfjLD+LvA
/0+83XjvRStFZYHY3B+gMhycYHfoSRBZyfnhG9RPb6RJLaSWHUuJqLCA089VGfvd
1FD4TE/3oycZMCrpqzQMy7GpXo7e9wOTNKrT2EyfFtcZe3Svot53IJAdc04WuT9C
17tSxJ8xgddGz9z3edLVGL8QT7Axm/K/3r7WyHZICZYa0DICCTSfETwkB04e32oj
OQ65cR/Qbzvun9/GDs/E3POcRr1bjktumjYWdjODZisYv2ygCtPy/38TfIrFBwdT
a0xL8JIPYYUqJQ/m3ISZTnIsa6VrnXeo3GmLQopGISCxpJuOMRxc/C5drOSQStXo
laUXT/mQI2LbzVn/mU5LCGRuHkfO2T0bNVxzDLGTOJwebmHjaILoDhgAxay0wAlh
x1GVUBJsa3pmyNXztuDIZoclpW50cINMX9j1JgaupCCSNvCkhs27KsgW40RuLWGU
n3jtzgQp8Zz0I3Wbu7CSjZCdafsgpK2yQEtLBrf9UOD6sVJamyguUPI3mwsW/84J
5cUDWkyqrEVMEotlCoc8UqUwJir/TO99j0mYqokRIpEFvpPeAUJU10eiQLpOwua+
5nKqj556mFmgXCO6SIS7zhkNo5UyB2efembizjn7VxLvokmLJvMpuux0Y5Wkr1Kt
+6FKXSxub+uqGuNaz/AIIU/C4UHU7lqPepwR46df3Y+014oJZo3tiE38xc2eJ23e
agDuKEUzLzZCy0F4z8pYpA==
`protect END_PROTECTED
