`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aUjyuBgpamKhL58BNYccPBqaygot70+keE6jIs1TOVgC
s7fu0PnTk/iWXiyyC8NfUbCDwCZiWni0BqY67C7Tj+BcCpegQ8NNQbEFR3/6R+Jp
IXioMNSOPJ44pWdCa+OP0uDAIIBwE8UyLSsLfbcD2ZGQ9LuiwFbtiB5m5kPFgAeK
MU4QnEu42ovGU9QDE4+OJWATRXCxUUJjxpF9OfpBMmpaVEGplFr1z1GNA/bmi0GM
b3Gdrym5mogxoL20dvhEcww/yAlfppLGlTb3KA/nLflA5qgfO3sSzMoYDnWSAwuo
WmHOyCul/4SlFRz2vmeB3ooBIi2F9HD5A6V9mLkU6qXziDoHZNJ59vsfr1ZYk9Ln
kMzLmNRjbP2LTQZ/r9tVBsInSsCu3s+cBVvTrMIXQbL8TzBk+wgCK6gNXx48XXkp
ri1Qniw9B96VsqmUptnTZY9Fmsv4ZNVYhCmnVpwP61xiwYJf9ETBYV4z6gMqHPwI
vDaCZzDH925iEVEwLJIKig==
`protect END_PROTECTED
