`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHlzU4W9/vYq7hoKaMXgQZ4JfAf+OjXMfwouIEUEWkGi
+rnk6fLqZth+i3u/sNu8vhN6px4yDOjAxuhwN8F35FfwE7t4tYJwUVlgStZ2/6Mo
E/LZT1MoOllcu+eDqnOR+pnJjMUlUajRp1NT4OrFiMxaf6i7J/1FzkqWxmh00kxl
SWOx54v416oyDlWa/IzgksFbfs4fbrf1ucBhu/tT0Zc2z6zghz02twZ7ngEhW8pw
`protect END_PROTECTED
