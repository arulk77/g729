`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDL8rvQ3FGvXRL3xQsYLV7/GpEQaC7L4HYw6ftGB/v+8
POiMv3yPBaJfDe3/+qKzrFUtvi3QaC7PQEfK4G0lAbp3cmMHQJVQI939W+R1eLIz
dG+EN7MKuZmNyuOSsFg1KEFi268YnXv8K5DW8Curqq0PHheYzHuHodIHT6DnfgSJ
rUHCsDFdHR+l2yAv06BEX1tcGhDVUQ+xdgPur64lEVw1RzxtELQL8koirMrmIwTf
K00OOpGCBS8FVlBz9RPKkDLA01sOBIdzli7M1S1Cjadpnqm6/iB0Nk1GQN8e7po3
r/xXmapFroHxpTve5ixi4lxtkNEUBs9OXuWKUzBgT4WkYVyJ5h41sQUt9PbTDkZO
wF71QnhE4nFjNwMGxtDSzD6wfyq4i2lR5YRPXeLGPUk/q2oNlAu0/FlWIdzN0v5t
hOj2Jk+RLGSznONTsUutTsRTnyzCREtFzQOhZZzEUyBlu3ggS3amMQg9EGy+tFj5
4xmG651/Ax3DpVnlqFSDwVjzaN19HPjxi1Dytjr9TxhqCmMcNHyflk/tIiKKmVDb
vX09rCx1itInKJ+i6qJGZg==
`protect END_PROTECTED
