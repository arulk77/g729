`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4w8a+SsIYuyjeLq4aaEfwnLhvx7WpqIBvbBsc4YIOLio
YR6ZJMGzBgDCvHmwRDGwjXBQxdZaNovM3Trkz778j0OuH+N4s5YsqaDdGij9ACWO
CMmqRCLoE0CPfYeoiJhC/kf4a4y9gpWYUpokE4dxiX4g1T11tZxzb4FnZEtDfwgX
5ObibAB2i0Hp3AA1BXFTfA+Uaw4UKCFsbrsNR2i0OWZyvYb4Npywdg+kNc7viJsL
g2ZeZ8tOJ4ZuUfxADENdg17ZYryhAi+OMv/aW2C72jrbLUXGIwsH0c8RDe+8A99x
6Sj8V8xtDUEH1PQGCoQH1A==
`protect END_PROTECTED
