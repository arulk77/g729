`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHwc4FVrx8f8tZVlBU9qcXRouwYAkVhBfaBNmtoeosEO
BshghfQmSB4VQZDhTVpfzXQvOY7HGhtStfwPE6CQB3oHeQcYSljKTYJREPMN5fzg
71AbCFSDoGq4jo3Un5Lox+8zfWZXYq0eE/8FLzTBKih/diD0Ddg3XwNVbN2ms2hC
FSetuPH9V2pcAl7KIHuZ+8Zj8fU1erMIDS5HPHtRGn41GxCCSF3NOAYKKEUmt/J4
`protect END_PROTECTED
