`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC2GZWOM+0Pel4+pJ5u+Wun2a++IMlfQ/IyJi2qEejC7
rzUDc3RrLw9Li9RKtYJBM2Sqaa/5dNnT4RklP0H9C8MyjuSxxiWWFigxrHYSbIVp
sSPlNgm7nL5lWk3NXulNWZQ5JPtyhDGsS51Xcxz5p7vTrBV3atg+Emplj3MDIylg
U6bJa/QAUfuPwuOUN573ZlmFgY9Yr8kJeGcXZ9wyDN8Ffh6ijU+QlWBgzPWfEMP7
NbHldxOfVBFO1b9MEMm8z0laceweQ3LWKx42yEPSTcKDnqLuxYHiYAh+9HuRdIB/
dVMw6lhklT6fm49bJkHYnPvbLmD2CjfF4Zfxa+jPTUFh0uyoRiHhtQttpLO/nRa1
xad06RWcEdlg6m0h90Uv53rDZr5gf53M45Q8YGJshSeknXnk14iTQ9krEyXDXN3p
a0c+SOGIjPH8xr1A652aiA/ROkJKLmmQ77staQtux8Wb30SwS+j1n2N/5MBMbJdM
U4rOajIwzr7M5aTVsdS25w==
`protect END_PROTECTED
