`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/nIjQvlXih4KQvwKiXxCITk9RCfPQ9TOZzse9sBmGzJ
rQW92CI6b5MDD/bfTSg4Q7ZFDR5h++WpHEyWoFjduoMuSwyg5+UV6jbJkGX962Zi
CeZLnfOaTRpZL8h6Pa0+gBaTkf5Jn+9ZbY+RiCEb/l0qR12jZV9w7rKWoOGzCI1S
OYj5LDkDJutBk1LWGLnYGR5jhBL6UfArz+3hiU64SekArQBur4iP5Wk3wbbBY226
lgocjclBFejK8TY1b+TlsjIlQ7ehf+ihs3ydeTDqlbfWXVlD9aJmbNO/S4xfyY9e
MP38aXkWj4MtLCUf+Z1tGWucBEALyMKqVI3iRy/l2Oo7fhqfPt+twheibDdMdPaT
KvHKWMRTc2uLtYFg6Iebdw==
`protect END_PROTECTED
