`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB1M7/AgkfG93JWOcGm9S8+NZVnCzqT8z3wu2+AS1Eaf
3AEskt9l+VAXM1NdsK1SRQNrGA6AiAzpQIy3jQIAPM45qYRRbb6muOGbKr9kzZVO
VLAnPJzbTG+AjO+Tpyf55n4Toi9ohmj07BPkkR/T31Hmq/r3QqBvNm98jiv263lB
myW4H332GUdlVLkx5Ghy33ibIBT00Iae5/TjMw7hxhTe3pRCNBruQE6/5D7CV6lB
5WEdfjpeFoRMK0aCjZ84lj0tUeKnb4s9jLlF44G4NGF1c596LMZCEXGhr61bYudp
xoZI2jD559CtLxXd1n5yK0bha/PlCJeudcOPyOjVnBONZCcbjlEsxgXIFy+AOe9o
`protect END_PROTECTED
