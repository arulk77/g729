`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45IbdW+I3npMndaEpKyrPVEXoLUJhYupicUoYFMIj0Md
T4kq8i+P+5LYrfa5MKN+gXRf8EuqMrauQiAwOiJHCx+3TDljxuC70/v1q2Ip+5f9
bPdbqieufFJ2tcnZmmPb7M1NyF8+McsKkZ9iStkov95PTXbs/g0xj2PcP4tyGCYI
V/ATKO6xdW6H2Anh3ZFgXvGliVGBETDllCtTCKsie6VxVeFjzVd+OVlN7mAvqwdN
1Gd7ssJGr0DeB4hTLNGOWMmiI1P0w0Xg90g+HOD+YY8=
`protect END_PROTECTED
