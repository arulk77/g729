`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM0XN3J1ISD4JFzXlSJ3pO4KWrq8sx9HZyQY4YRiOE1t
hW9+wTykhjy5y/8iMSF8cjsLK0I8pAfo9Z8wazqch8E1vT0pdpW51hcWXMy1F8yV
ZcUqYl3FNPa2us9Rj+peL6P8gs36gJF26JljRI2wrgc+h0ZALKW/+2RpnYhCy2i+
`protect END_PROTECTED
