`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/QBVX3ZGTYguXpu5Taw0R4cXaUt/cFaoioqbkz4qDnN2
zOFDXzk7QZ12a0RVH3r9piffaJ+YHmoiVlzGvQBLpZKkhmnrzqTZF01u5EtMa629
O6qm+gQ3T/5dfpH9YfASW/dxadAWDmihfY6EMb31c7FKu99d8ItfMic1FkZGmEjc
oyWKBUIlhCXZIAzFDyJ1zEZetSf146WiFOSB+rMDK2169KohjN6uXxa8RwxuJs7A
v8qhx7yYgzW6kAHPWO/CWvQAHlS9wpNW8ZpI7pTQ0yJWV57HsEJ03PmJTnt/39wh
jEg7mXzoLf9BYB6x2gs8G1SPNIcmmMrac0sCX4QezrZGwoDTqjXUq9XAYaUFWKem
ZXblYNrOZa9c1zu5Azd2vjXIfGNXw8FHbkTtxwpVTbvekB5fJtHibNYrY7Bl6We9
a+PqRBFXSDWChOdmvD/lVW1mfAuKfSumteWxwpwN804=
`protect END_PROTECTED
