`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAVlm07DSGRUyulpMZ37x0dvN+rxt4zVHqEpXf/XvG77r
MH63u0A8vyMWlqc795KTR55PXkgJMYi14nJvTT5d+UzzK1LX+caMahEfLp0IgyN0
kVhGo/bGdE2q25slPSnA1O1+ecN8Ugj7ROgYZg2HMbv2vHkBb63lsSPybxpRvFu+
/dIiVS9HtM4JUX9nL7LVza1apciNfPyNI5BvGBYXtkUxpeXXLi8lGIdDQ2k4j3bA
l10ixuPwLsqJDQ+PbgtWWctndcoLqo8Cw0DmkGpfbg91LPZZxqbMOubl4MefWtDL
mJOd9kZ09KjNvZTcDjia/p1u8ZTIYhCUGOTW//G8Uu1nt2pWK62Vr2TuCbuhFGT5
X2rwozoFxQqGFXPNynuiS/seI5/+y7juv83wD031ccTgc7MB5zaZ3LHHmXTGGG3k
mrkouoW5dUpoF0BorMFJTyFi12lTR05My42bMy3dx9cwFHyUHpCYR/5sOFvQgonm
uUMVX1aP9oBIbJvl0Air4REDGgmoQy0mCBjI/WIhTWOzrqc5Tkz4PoAkUEyZvquf
APiK2VCUaihxRo5N9aFqAOEZTIrETRO3EBjW5eiQNtlo6K7VBxwPzTGb92PDTtV3
SbA0YfcdqBsQGZw4zHNwZptOfHf1uxphtcc3yc16AigdqpyXj4iw5neyyF4hbARC
fpoxN7JV41rxU7dWJ8rmt4UFT4ZvqIhNwF1Ba/Jd5xe8qYyNqYJ2zBpzPHtq3G0Y
pXaPyJPgOyCS9tIslWUVYBhMyJWT75q3a5P0dfwUkjiBjiMSDApwKA4mXVTsfapU
M8TIffncHKrWSenEnagRBXMQ7JJX9Q+Zm4y19pVZuIiu2LHlt62hAB2YZ9pvOP7/
nI+i3OP1aygr4MWON+aowKMzt6tvEGvbZNeWpQiyq3V7brVa59WwHSu7oBEdb7KZ
mK4PubmHLpEW447+4UJOQN4PyhrxJc0dQ6I9Mc0bJVkIokLFCh5qN7oqMqSCIuKO
6998gBVdAjRUzz/WCwmAioeJwK2HkVV8DZzAkPYbqRin+/J4dshnaCYlQcUmJKmL
jD5c6Kwy2v4nw0PmrA30jzHyIlfB0MKqkXsJx+KCyuy0S8JRRENwddsAVM0pXLcR
keqxlfZ3iThWPlxt/9AYGJJft//PMwUwm9Rlf/m2g4QIVDEmD2TpGTlngrgHAv1B
AGfg8/Ki5pbWZwZxA4t+Kw==
`protect END_PROTECTED
