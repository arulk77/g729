`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
spj5cbr6oJS8rhdiClItU7D18BOwmYaXGjYTpgHaE0hROzYIMEG/0B6gROMtbCe6
YYY2k7/HPo49gfOyQAfTPKe80SdBJCMRgLEJV+G7hCwzvDuG4MtrFFJtvLxHzKzC
qdupZj8A8Ws1iGMTOJ8IsohmXvNidktv6RjwlRytxQluEv76BWyazmpRQ6a9CbD/
6nRXXMPLE9QcD/5b59kKVMOfsAJHzSjqCnD6YiTwmlBweMhxPVeqrJbDMu/d4Vc7
yOfLZL1rloR+x1suDFajXh88Nw2u9+T1o0rB7n5nX8M=
`protect END_PROTECTED
