`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNVxEJ4ZOF64oIg2w/cSzfVBkB52450nK9ExGMvGg4iv
W3H1INqq5AwJ9m5VLM+jyG9cjI3sd9SItU9W4fBFZWmKMTDwJXgPnkmY/8PvW0Ri
2Kbqi9fFArXGG8u8o6YqWxeZVzFFbJTxU+dnYEfzCYM+tnWiee2yibr7PSdDgL/P
Yu+edCSiFGeHJQzT0k2ZSvtoARtGAz4GYT6CKrl2Wl4c0nrYWyKsDo+FnRUOUcTA
qDJbJC8lTmFBJzLzXQrLmXYr4Z5knHpkiLDRkiqFppLSLwT0EsDgwswKoDoBTMHO
aafhs0D07j9Ay061g5dcZvkrya+qIi3Obwqsg285pF/aEcNedq4aPf+VcYItDanh
+JPLHe9QfYyZXBzHmZZObA5L1kNx+wqGjMOBKA0rw2BX7m88RPbj+aT+nEebf8GT
a0wFCAdcaUQ9R9AXK2kgv+PhdGQULYdCRxE/jCiT4BK1GtHigrrJrDH9chO10egu
8vxOAo5In40gunIx+SUqAw+CiKyVY+CXK2NLOOeU1mZGej0daQ3EpzVG0b7c/Kso
pdAIvb28umPhcJA9tUMu5HUTl4vAoWMosXK/TpWizaviOtRG2i8a5yZvKsibAcIu
0uutDtxyrrmf9hTms2UkvNcTKiFIEHcGTSe2+b0kU11sbU17vyiDB5oXdgQtY8lY
eEhFo6WfBcGk31jszNSz5c4JWyrD6p5q/RyNWR8CI/K1aIfgPfQmXbWkwlUma8dB
V2vLBah23OoMkRWMdZ8am36dp8W71WS32P3Rac4+aCd7wm3Ura7K7XSMsrMYo9sN
din6koRCjv3vhLKDLG9axC1JCZ2Y7H02zmSKLdtBLKFtZtK9X+ACPO6EqXy1nG0e
bwTvqCGB0zduPbMPs+NeEPFcIwfjOxOupzGzl0plIkNyjFumYTn6iHopCXzEtvWp
Nkwr4bUJg3Bx5D3+REDNYHAJ/fkPJ5/6CQvgpREzSz6h1ms5rn76cO7iX35P+wcS
X27l1S6xyDfk5LEj4tKWy4p6gCUQeN31oB7CEpiCbMHGPYpXlvD2dFE3n3eWAF6N
1dWLzFV2y2Ihg0RAjqNKcikYEPTmGgoGq6oCS4VjDfzeXr3RNcc6nNdnnf9WHIbj
lDtJe1ho8VkjFegFFG6t3d0fLu6jgq1zB8X4X3fRvM5dZ6jEv0Oi32iClfBH6xZB
H/Dlnvl4I6VRv6Vyr+renHjiVrnfmKfcCHDL18YjgEf1+VK1Ui9mvlvspiN0qe13
h9hLCayuSW+PfV1FzJKGJqh2NeEGp3vF4tYuNQB4ubLn/HFVhLiBRN654LJRXFc0
XCi14pYfexxcX90JXdBN5+mABSUBzgJTVj7RgplFYz0DCA1PiRqzGRaJ2MgHzC7v
HDr1tUy0JWeYuXNjsQAuDcgaWGAXCm07st+9kr23YHnRn8Tiu7+7Zs3BJ0/kSiMP
VUCanQpB+wm4HO0r9YvotprmyWGUNa25apTks+Vs0m5KkUlILIYtadwMExrzEssE
ZnpXEQqTuQlRkbdEilDQIS678MiF3N6fu4reNoX7JnB4Y+wd0di7D63WgnjDfoFK
0hhP7OfXlnd+lWmL6Q4/oEkynEIVwgctWoyZA1RCjwOEwi3s/AvNzM2vVLpFRlqz
bQV+2cwQjoZSDePNVYnEn9wRGFPW8QWi0OHPH4IWx1w1/fc8qI35lY/7wXyKncJ+
Q+vD0HBEctcfcsMtMF9Zs4uvHyoiD3KNAXz+LRgVpNfEq/pZJhqqccAXh9rJJ24G
1f0903KfCwL2OgeWLdiqFlNhKVl+Vzzpt5ulm17qlTwVuK88RSc4QrCE0M0jHTvw
h3ZRHGPxBoB5KDku29WKAen9ZZR1DFp1j4mlaW6sw7GMe/Yf0x4WJcASGG+xR0t8
fwFzyrlXCcZHic+jViaO6ZAtpzGw/vAChvXcTim3cx72srKqHLsb1bKIeUFU+6Nd
kVDu1gyTZmg93j3Aca0l4++gN1loC/box/yJ5S2PBe2I41J1p3NYsD7gtJMEyrFu
4PRvSqE7KKcx/cQoxpenb9pW251VjuH8VViOGgxA1A76N1+KShCNKm9Fl8PTgGIO
uGNdciT6+XriUrzzwEbitFa7lfPYiXh9MbmG/FWoubFmdsnwPloAQIhNHR5GFX4v
E70h1jzbTUkMc5Bs0vG2rvRM7xw+NJUqnJUPvMyPOwEMvF76PfTVdxruStFhP3N1
TirmYtxynHMBH7F0nJJVRv/2lb71VAFD2PfZo4QvcCCvMBY4groHhK3zOgi0/2S5
03vhs4lylWu5S16+qfTds4XOu/BUJ/23x7taHuzZGowIgGq2Ik/01vjWxINcj4iy
PC0tqp0krBnZDWHI19cp2WJcNVW9DNhqwP70uSKejvrcJhqrzyCmYCZZW77ewPtv
0HSzWjoBlVqnFcHGg0aGvpYJahvDoS25+RF7miQ2EARpeh7cKYkhXqG1GvXbIn0h
t6s6LLpWnSy2qgU0J4A4ZkJi5DrA6GLze2rbCz3LxgoXS7IotoeX0bl65sqISlk9
Z+INer2qLboPP0DIQblVqNWtTqpurKovNTWKASNylHxA7ALFoDSDuZWoJ1sWRUAp
NRwWTGHOp7EXaDqDnNpRY47UFYJXfKdJ8bkIixpSfKdEF+fztvckYtKfT+1UyDVP
xdSxuIa1/uuUG8FcQMXQHqsQyUQ6tBaMiRcNVx1FPNUU/nvhQG94r1zo6BYYt1Ln
8c/v2ILK8QdE4L0DkqcGFuK9nPCsVbtuLdDkUbxKzZku8d2QSH6nFvb1DEYuWBSk
jclNCnhS1TEPdR8LVdhHNDiaR2pAcRdqB7zEtcoW36LCohxF4RBT8MiCI+DA420G
WjZYzii/3J3BvNOw4vM0jCjpbo9osykEhY7J0vApbAMZxVmlTrFpgh3okH1P8xGb
8r7oEHtmmq7n3BKqj3aH0A==
`protect END_PROTECTED
