`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+yuK1d2NT5NU1FEcMoBs6CZ9G+9w8yWVQdyxn9N7AKj
Aan3gj2IzhJqr0F+emBIiW3h5n2umN6n4w+Hj7R07cAWYJV0rGCac8OvrYjvQYu+
Se1Tc+EPGrI8xXvDZ7xy3DdrQfbD2nfYcaSgfEfRuqWuWC7+CRaXcy17VAuHOlWs
25iYPrd9t1vAxVzqgaNKG24dGF3Kpu76KloTGB9jjrg=
`protect END_PROTECTED
