`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/MY+69gJhOa4DAwnq78jVJ8YuZUMmuz6NGz3jIOUI0+
7HchsP2ERoA7GJJ7D1UNhnZxEnzoITTkN5wq7a7hfm9MvF/T8voYxW176T9K/Saw
JQa07gwBsUB/yOprACh5unDYvKR3IGgQNFqrwm2VbxcyiEk80DN2en3p1GYpDah2
PrvZA7RS1T/dZY0NK2U8IZz3y7UromTUOgRy2wy0DdnbzRvdTu14rLN7qgyWwL8M
nnQiv3O3vGmj8Dhw9O0jjbg9E4/UquXqlfLv2kxj/itUqRn3fFbBAsB9Pw4sp5kc
+II2FB5IM0eQ7oqcLHdKtJkLBA0ckW+PujTXfFknknFy+bk1g/F1qL9gJXef6mgV
zph1+D32y5b1h+xIbXiVlw==
`protect END_PROTECTED
