`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Rj142sNDO1F/EvC9ghDRuGXg5HR5AwpmfQM9xa6UrEphtY85oLbVzA6JiBhGA5pP
C7aNVqDOLf7YKCHbG4QSCNhoptQAGGhz4KVL5HQZxzT2v+NcQW5/8iyOEJmbftNa
aAMYSktkAk+tLSeNzcdzXhmyCpO4dM5k5T3XYHTuOd3tf+ryPbHPWAZbHkjHVvNa
FgvfkpLAHso/OEyEgMvMOuI/17BN/D5EL3IyuGD2u8p/9QXFIahMBzpX6wChnLdN
aEXLIS+gn3Cqq0Eu5H9NMt9z1gIPy9j0PGZvDfU2e0ttefAEnlQfg4SbQArE70Ms
/KXgxjW90eYBoCY5uCp2FzwfQEQxTZIl24+yQbxufUuvsdJd8Cj9EivXjm6+NAVb
23QFgZiT7E5cB4hl5PfWRgOds9BxybvHar0bC43I2iqVatkzxFiIbqM+F3Rh7vjs
CBF9Kil+2ilnODLtJvIPM5Ytm3J16PMoQI92a96EYWKXf85liZe1OU0a9nz6SW26
myc9AT8m9rTHr5xg/jQAN7KwB5qs2fXliEt6pe/N6hqqFXQezkU6nJVoQFNdI0/N
96ArSkzcZVBEwfVBo8Xbm4i5nGbw5fvBHPbSX+lHRFzAr7v5+cKp4Hg13WmN4QRq
C3KRkn+yynuCdeuaERs167x8d85JRqwPvyBH+77bq0dOsILSlVTC489Dmx12QG3n
uwalLGo7XckpxREsd7UOYCYt0WU8dne46/cAR/wLWThsuNeWpB3e17GZTRTjuHIb
aSsBwQbnNUt63+yj9zkgmm+6j60S74ZNnqypOaewifsyM8YMfxU6FDgnjUmOBzdm
bgt7GySWHjfvUm533bEUwEwU7i+4CyLGe5n+A2L7tTaMpGh2u6OMqnvnDoPaZFPM
YPShVpW/RSnnrGCt4aiX+h6VOdg5KrdyZL1RVC96KyuQswqgsVAsg8nRjL/47NDu
wO2XN0CR1vp8ZcAODidriMpxrGl+tRZ94iTx7wHAWk3M44Q6bW5ap/JVkwYiBRxT
ik8txSEw00m8rvWJSnbVu14GPFKJcRftsAYZsUjoY+DTGwDw0TadmtlD5hIwK657
Uhv5e2AES8JHQyghIJnsnPGYa3CsiIGVqAEfOVRtwqylUP9u71QkkTJisoAp+gdA
by9s2+65KzCMFIEDL1DvAgGtNWkoN724l9ejM9RAaJC616yvITUwWN/J3o7zA7yg
S8mBcFV9YCsJ9ry0IEvVsrAlIiHBVRWg1pIxgYmfSeMsGB+G7sbXWL5QyUkNlI7C
JaeUcRFNd6ALbgOlpl3T00CgMUPHU3FY6r0ChFxKqwoueR4+PgZa5gMaIuLOXEAy
nV37h0U1lSKF2elNlCg1qL6cJvYQwzDLgzB8adNadKDxJSFomBhYus95/24HTLdg
CXynUQcHkW+YvpYAq2kk3Z18+APPWF6HmQOj/RYAIaPhmy8esUY92ZFIjx1mOUB8
UMUeURkYCSd45nW1XneLuJ4vIziKpIdtsvP12/S0wPVUnKiJB5irobGEbyMP3Ytr
eT1KfsWJqNoM9c/oQghlzwSE8tFvShYJrC96b3jXuzNFzvdtOw0Iet29/SqbJ68U
r/C64Usv215x2b8XTG1TiV1Rr6gfR/aOIAPDz607VbdlOhxEs0h5uOcKWQN28ETJ
0zh5Fn7f9yRu5doIY7gCwatBUVMmT3j1D2RTfybacSAYGZMkIEmfpRZK4CpoKwK5
/VRmCEdffvewT7s58CnDkn7qWrmi8aJtsf5Bkzfap9UALXcKTmXYIN+VGFgpQHdr
7ZH+yYq5DtUhEnUD5tA4qJkKibn8kE9Yl/34/AXY+tW9tSBD7e7Z2kdIw8BB+Z+A
SkBYN2xIDgo8LzquYPc9HkuXBamJ40Xr696z5XqP2CEPRMC+xHKWOijDxSJWlBZ+
qbd3/yKQHb9gUu9VLrCgbV3/BqQG+A8B0cG4sSpv0sCDASl5e6W+gST0IbhjtHeZ
edVa/JvkhGEx4mCfmHIzIhav0x0BvmoR0KgHoRKFe2AWs06+ihbRHDQuWX+HMHfL
AS44a63yoThfru4mTwxzwexCYj7KXIal5I2PrEy1+d54YAP4GkghvDKVDWyC1NpG
o22Ld4fW/nUmgyYjZhYs2aZPHGGem1kMba0uJthFZO0Vhe2nxIOGTQvDeNTL2Gbo
cHN0MMEUBkqyEc138xr/QQ8LDHVmTjLqgOtXF/hzDG7yyDfHqmg09rx615OVdRs3
OjfCplh7QMNDYR0K3AdwhrIo5Xh2l0AYeGyhSc1Fh6XaiJ2hSUoi56K55AADFHOe
8Ygrjvz3Fj3IgtYHis/Bsh7EFS2E12bdRhkIWx9EqghwPGGbiPlTU37r4SRc3aLJ
XhfV2ZgZHK2fTWeXMBp+Ep/ZMeIvwF6GzJitvTOFPSDa3h6Avx3BdDyi/k3NA335
d/4n42mg4Bhqdpk9PM018xUcNdhrYygOlOTvbJhb9tdBoNKXerZ4XCKobwmjSvut
vZJOmP5Yg3nPbPIz5qSwvf0o8Y+9qrmVLsS2N+jSgW1iJYa8imocp6yLLZkuJZiC
EUV6lwZfOCl9RVWuhK3Zn4pvTHD5bj6NJMg0uAYULcnxIcmnR7ZIFwclUcp+mw2l
jF88cdFY72oMxYkNFoXWR/KX3BKaOJvR4Fx5yn25y/MdfKS3w5IlaTT1lRsaBCjv
LhySY0+b/OcQ/K6ARI4DvTY1SAsLVD5UD4MJ0wAE0ew/7lzFfSpTrZkjhBesCV6L
Iqcpi7QWzymHLZ8xNqkb+5amVFSPqBzoykBzIMdSfW0dfKwcCrNgZoMgeF8TdiVc
3kCNO5jXeCv9Ayplda/kMPd2WWsZ0lEMnj1OsadUpDC8VdehmUrIfOdJ+KTQbhoq
q89CDCCltzx0++DVt3aUUgU9pIDfJllapgvxNmLT9Xc44jm++4qjh3Qu+/7z08Wg
vbGCGid+f5px12LlXDtQBkA0Yiw5NfL6qJxkYzSnVI88RhZuK5XWo/ayE1HrkMm7
auPVKmLQr/wgEFXpX5DbgFtUHWugxx56PYh+Z7hzB/wTuwsibCBjYSRFHKHnaYVz
3pAcPv9VN3R8ATR95CaxwOPQXNMQKOF+5/cWzBVyhQEddslA/W39rV39kHElTRHK
NIaeaJir3aR7dNb/zi34jbGXUqpIGd0FEBLCJDi5NQy08tHymlCmxO9HPu/F5WyC
WGbLHEmo1WKdhuZ5QDV/5uogoB6zLutqobDWZgGybReW7fjxn4FcF1E/kZQBKOdB
1OsEC101NwAFrnIHgbQxbdkLdp/wuuPJgiTixrrZFygKVzc29h0Ogtn7TFQcY5a5
uiqX1weBM3tZ+hd/ohnOJRPxEX675ZHu48TaELFhi50nJiUXyWsSPARpkbkjla3g
2hEYvaO3gT1FxJcvnP9S/QO1MdX2cSReN2vWYb4hr9ht6Ku7WaG+oHmLwBOZ5amG
5qwtGceI5Tts02Kpz395Wy1jlqbIv9TCypiHdgWuWr4C+OhuepqJjK708vlIVuTq
D42GfhuDeHTDlXoARv00lR++U7GVeySTDNSQacAcFMqGZtud9zfBekUadZbytZSJ
ZboB2yyOFr1/2NuqQ2B0FBTz4qv+0DMqimZMZsRcvJEnXd3tOOd/dtK3tsByQkwJ
2Wt/WDqv2OMn1cMFpZdSq2Pkx2SOv25C29svmgFTIVl+k3CFYdmbWriv7VH13H3K
nV4Cce5hSfEpV1xxsa4pONwPHU/TwGCTOaVdAtHtTDQb6TQW0IMc5iNfUioSwBBr
xMREx1UdWq0Bwrdp1UiazDivIhAuLEZSxD8vQQGhHBDPdNI08N1K/N7EgtCkPzlj
LcOKVzwaCp2TKSdIHMxFnhF6Ih3pjYYigb0ZlCdbkN4fkqV3+5DGQEEdtm7lTSgU
pKxOKKgXIfYK6Mwb2HLHgt4c9728pRvmiKMAJYjK54iI0r/0XqZvVn1q+EVLyuIk
h+ZfWqFY7PXp2OlufN7hj7WHDbyb6H3Kj71kFobWCw9umVgo1+9jeKXujyL2J4dQ
4AuoDR/VcPvglmPfM9EjpwlBmbsX/Srr4GEaRJaDxVcC1nFxE8D385dgTAdMn130
8wG8AHrp3fqQiBtJ7ZFVT9xN1Oh0PwTB3Gr3pvAW0mInCykHjFfZgEr2cM/3vLsc
uIcXh80XruRFuF4fpkKI8nCePHM9HBJbIVqh/H8VdF8wtA62Oiq5gFB3VNVGrYho
2umUyfxpuvrVMxnRx9MhrjDyI1CsXWsWa2WfgERMV9Y5ZHLPSizq3U8/1NC+9OSv
EDpTZgyWUKSqmq1RXpVv4dLW9ExWFZGnVVZ11NN5AD4YCfhZhI+uBhZ8wBUDXaEL
uWpHVhrOtp28onkZzgjp/zqigFJfkUzWOx+jB7o2DuYqe9oMQpJnjbWLTkPjUZpR
jrJCUHYE1KOieQ7KkA5iqg==
`protect END_PROTECTED
