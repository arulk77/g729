`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1ad5wy16B/1WleGVjopfXhPs7aKSBQyJAQ2CAGg/87bmZ
BZxjP5PQxvIolE+U4hNtletJIuMuzwJd14hJ1SJDpPiQEl+pD1zwqtIFb/Lg6fp/
H4gocZZ6Msazs93sNzhOhYkMFTjNomBtRf126M9xfQ+6dn+Xig0DMqA74cdO+xvH
/s88I8SuWIOklQDuMrtQhsY3a4bLIEuiuQJ/kbltAMh77VLc8a0CSr3TjUvX6N2a
w1Db3sfj6YgyEfvRpwo0VXbdXpEtzCfCVmsbMoAqZ8zGavKDmiZvzTphAllgiL9N
nsw5BW+Glj2a04M23RAVrhHdZeNhM5fCMIGhX1c+K6FiRbkvcraTHdOBuJKpxxZ1
zdTek4yuFD3A1cObLFd3EAfKYBfknGj/Gw4HqEbi504=
`protect END_PROTECTED
