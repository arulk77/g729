`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBk8Oc4UDV2/5nlxuTR0RPu+WtmYEMXGskfcR3X8x9fp
WgJbezlR8gaBNrLr35af97DWAgzUxUQvP+div5l38sWLhMVwkquJJBQg7i3ebjsB
aj3tVqVcAW1+0KHtyRRZB7/tB7vzo1tpWnpqsMloKyZsuHVmDt5HvT6a5mAhjhAJ
`protect END_PROTECTED
