`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEtFC3ntBfQqiGX3nqUHPaHHFXzJJtnQbb0AEwyu+RQU
dpfYCo7wpqMqPcdhkPd6LEp+hHJgtj3BlEdMiQ+ZSnvWQNcwCbKGUSRnmZxCnc61
o6ECSA+44yWhnXjrC3lr9ALSPZXZ5SxdE9IPK9R5T7prLuzpV/L66Bk5Q9k7+i/f
nmWJJBUSg7tgk2Q7LWOhU4hpLn+K2/A1Z0/grw6PUuOAUdQI4wTyzgSfgmAh8zRI
/VtdgBoEH12lfQ5fw01rUVOO0REV9hYpCODwBXmKvEhX3zSNF+F5St1pdbpKiITZ
oEAC5aQHrqFuOHFs25vNCjg4e5Lxal4YaHxX/ApBesJCWW11ebT2Pc9REUb0enJV
`protect END_PROTECTED
