`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAXxZNlk/x11kpfOsWbgldij35nFWL1bggMTcabWTYPdA
OAU8Gr6axUDvmGxHPdLl9zM+zd1wi+QRx1hEsprI+Ji8TJVQqh4+260MDQtso2yg
d+sEEQeDniDFeo1lvufbMArFR8YepnsyQKHYM8p44eX3FZPDZFTqVoYCa1uqlLed
3BnW2grt4I+28eSHds5VLdOPfVx+vHYlIGDVWu6XQ1m04s+yvwUM3h04sEhxtHIl
6Gu3A1qk+KTP3+hw7IvRhpxrTUtltKaoFYc5jOd58dJ1ryfl9rKm4fYsLw9x16cs
6qNRt5yaZHiHzWeAxU2LxEdHnYnSKY+3QaxOKSDrWq70NTzby0a0ra8RUlxtzWKl
yxcUZfTUG+ueTk4aQTfjLnAkZxdFwg/ikWsFExOWot8sH01qYyR55NXt6HMx3tY6
JfO7DjlkiBYr/iZtcvvaeGqrXp0qKP//KK4uL1h6QEXYVBfsn4At972wfU/k8+o7
LAEhzFg6xl61m7Ch1JTNzxKG5ZA18BzY36ocfh00fS6hFaRHUZjjIpqx7n0d2YPM
MPdw4uMLa3IpExKJhpBSxER8FzDPVOW2yvCz89rWcx3QeT8hsUt6DTo62M7bKvx0
xaCK95otASXVHhXnnCYUod6kccfE32CPcQN2X7kMu4uijARDPyCJj5qPhKZK9RAa
8P7MV2uxhzeqEBpqVEaJLaCERxYZwOtj6Nc7vnJv2pt/eM+UJdEX5YlecA0dJPR0
SauPY3m6PRwPPfS9CK6ugZzvq4B7RY1an0P130jvY/KHTjkKQB5mMvwPF2R7SMWL
lswBPCD7S3lQ1trCFuY2KQtk7N6oC2B6gymsPkLl0/NoZ1Obj2hByt9gPPoYilKg
EGlYSzefx3eswbXSZePkHIvP/CDZl6dOhGVOc7QaHcA5uDFfx52wjSr0Ne/HygeM
zp+PKTVLcQESBO9P878sMeWr6SMnnudjVzgGmrKVIHfKD7DbcJbm0mFcYmy3glaL
9BhW9fY0O2xKkBzcAKMG1sOYJXBaU3KjUWMiW0WxB1+OHhupoGRCPCh5PnZ2oAsP
uute7o/mfN+yE1mmZ3faLOdqCHIHBKP7+oOB47MpxxN3jDzjhx8uTJUiCgjKiDda
xvnL8sUkS0lFGaDgywKc4orIylW18009isOYJnuqAopXekGW4WOACGUQ1wKkVPYg
PFj0hqNJPZuC798k5evqCPejnCIzOvblIdslPg/7JSfj1qz9WEtwJ5UNNGX04TSO
PS2vyKoA+/8saGOwGxB/E39nRMURiIOC0sfuwxkANKWobQvh2g8TNvin6OwdvxEC
bOcO+Hf/ZV1Wk0PFBwV7E84rSm0HoP1p50cHo3BHPCRHsMqoXOD3mJSzBbxzTYHf
1Mqkkz+X3OP1Vq/FHBPMHOHbRD3Cu2a01Gun/xRtbrtBqrRBV8PiMQA7Pf6Jg1Ek
DVye6fQ3zGyBP+J8oDgM1Po+5cs5r3JDe8FzrwarORmobvR/HPmpgf25fKWOim4V
DDLE/2Gsx5RdcVNLRWfHQJykXOCAK4lgjX4B+NXk0jxNbVZy6xgDIe/XEXovA2hv
mU7apyvr/MoPJTy+WcjkrLG/Rr1j0Wg/3lv9FNf0SFAUs/KBUvBoSai5EHBfjlnz
KTwLB/jGXc4njwojzAl/RQr+nemeOFIZLITYtiEMo/uBrblUGUTtddDzePefU7cY
OWgn2PhZc0HsQ2uLmWQjuzNa/RyksXMey2TwR5Rq9iF21ERykDZtsBQPQwnIP2RJ
+cx+3hK1R4JriTEKOpy4krSJqqcDWOCvC55Wt7hvQ5md738oJ3ApZLdTLLgWp8Ke
4evPwpkpflDwO3sllzyBy77CjTKzXdrEhrzjg5IpdpXvZVq3gMZo5NIOCRiepx7X
rCi3pi7ji3NfElUiQ21Tan5wq8RSONL2yM2M8ZiNcRzZhGLT8Cl+ORDnvWmE8I/a
vUOQcVdVdS+EHsMV6cXlHoMxYCurSpjpruMpqb1eyFmuuDn9D2kW78SlGLfAS7lU
tyn7ibV3E5U2vxA0bODua5FalfkAVHCsm2ecHazyyzl2oxKWvZMhBTPy5dWc21XZ
TFEGKAu7gGTnsPiTLwuIbKrtMY2faV3VYMxDvYcDPofI2LJL96PFp8wEpNl8Sgwx
EoPLm0NNoledJLU/U8rPjaJv6j/4jImS9Lry3zEObNCIzexNpwM1yU5cEmHlqVmP
53uh//T0zqU+1PocpZXrSglJmQSU6ip2V8i2Qpbou8pbV/xj+82r9VNFB6Bpai20
WROpEI0i1kqOlR/WSPnmBvGDhMUHvVgvd+TVetZu6s+RUdfx3GSosMWM+nt1uGbn
G6gybW4Kdk5LiqK7MlX6onRBQxpR8ir89UTiJX56/X1RjdRDZR6Pr/IWMEYzrPVS
7ToZyht0UPl2PX1AE1Qyl7pIO/Rm+N0liESASJ8iY1BfVYDPVsV1wfkA2H1hcSnO
X+EAKTIXPESTH2K4g9gQD0y/U0oYIFKW2rO67f6P/PHTG3Up4ulWZqkYNDXqiHrW
o8mGL8MKpgN6+2VKw8S0IZzTcr0yI+435cZ+AJQiGOsJEU/ZBFmH4fEdno2Ueajp
eDo1zKdcLx/m+mnFnOaKlv9KrO4wCdZlISw/8Jn7cPafP9kRmCdyXPc6n2LfJHVN
yh7+RvzHZnOUZ0aFdnwDZQ9HOpR5W8RVEK/Yr+SOHpw6pAUrus3yIDw6aS5ASN2G
cd/f4Jo4NBCDkNoCNs47EXiiIdxffxD7pdznpF1XvxuWL9kn7esmye8RorPwqXN2
92gcqOsc2INbfvXvCVBw0PVRChhvLQA+k10Ngd9kuoIV2Wzjnsz597+I/Jze35BC
ODyeR0vNasM70SsNcgERaYF+Ru6oV0vVOfe9Qvnowqdodd2E42V51GeydOjdcdh4
8ltpAbTeIEcd4tQYInfgTg8jOhWYjNKRJg4PCjw/76LYF6VFHGcwUuOC/wmrnJBb
7UkQnJ1mwl9CfR0VVvRPVep/L5WBuN9zvEVcjJQpjtSLIA65XQJFemajYdX7Zshj
cwDVQ1iFnb++ECYDdyf8rC+S4GQHrSCXm3GxFiRw8sIAWbZcHe1+tIhwo3sK8h3C
DT8dn3fIfPNlcQmV9bcX1twwRDNS1vWjSxOrThdbZyfWdXh4FcyLKQ57NmeNFpc/
WoegKD0tIp1v52UK+UHNUsqgR5TK78RuVgXH2H1uwAxHZyen3hkQwS2oXbYhHKpr
a08GCi+nVV+xHKgDVvO7JFAlkBFo1VF0Ix1I4xxzuIJc6fdOmcF5gzI6U6I6hhJv
w0GzbgOCpdhNCOXrJQX+bbH7027PeSw+0uGsP2sxbfX2FiLiYBXTy0EcRQw5w9Op
RB9lXc/cYjjNusQGwlMoUITGQ0z3z3JK/w5jhLyNbVdupzeuV2xHpeTm2SQkyx5S
0KJkyvh8d/9naepic+Xt+jmzQ2RGPtmmtayKXOF7kYb0X+NxDHCioxtcd6Nal/24
v/V7iYzc3phsRz1I2osF7Tfcol7vk5/9MyNwR0aTSyYypQfL85uyZ/sYFqx0v+Lz
`protect END_PROTECTED
