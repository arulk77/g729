`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4y0tVr3+mhKeHaGIAWnfe5JwAQF9Zz3/w2Lh5dPxWsjb
SdxuIyTYo2z1zu/0Hw1DTAJ6q+ybwnBha6tGgP9IGBOMczPK3+9QvHdT46mqkXHh
R5Rjk9aj/pCc728DpIIfqJrYgJuFwPrW7HS4MrWj0II90Gli8ITuoAeC2rAI2Jks
6iMYQ/Pdw26paQVGnKbu0d7pD17Mgg3h5RxTlXwwUZ9PRmVNZVVHdrIZuyZhSpIY
NTAvSJAtbCAuBnLXtrBx8GH7KrSamICh97Q2NyfqCy/wqUPYmoE9iaa2aKfjiZzR
TH4opMyrQ7l6AA7g67OVqg==
`protect END_PROTECTED
