`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Eogy+zHDzNL0XXQvxbkIF5BH06tpU0ViIr3iWFRIOTrCBGagLfGG84tE1qg6G1fq
P2SJkjDC4BjnK7miJq6wBKoXi73fVOTFkVPGjXn3cNpBXN5qHF0At5LQSE1QxzLL
Adnn3m99EArKBUTSXtXlsSlJd7+uCodj2fHVgIku6YWxenVp/CrYDNHxETHC/zRQ
Xr4jpUz7ZeBOkdbw5Uf55x8D+MpQtcU18XnxMPd+Yb4BWwDhFfwBPJP4KmNhqGnJ
Tud7YwQaqbLSH4hshXtBphZDiKleDFlWUmNtCt89uDqSakiUWAV3fx9KSDuZGj/S
aFsBeQSr8gdRESOme3G0dA==
`protect END_PROTECTED
