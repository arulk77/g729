`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
l/mkjosXUBshoJR46TE53nqHwBEnqDVMNyYRT0+iBILOdfBck5L7h+cSgKI7iMCv
pg9KSfSuQX8oGj4bZIDML4tT67NXoieD6nVH5nlatsTQ6OdbofBvI819JSNSlFn8
Khq6+L+LgJ11T/8Z5Oo0YKU+WgFcN4Jeqe3vpVWTVLKUxiGLr1Ch1oQW6bVL/hBJ
Ffit0/sc8HV1MSQjgZDLQSnNDjibvwFe7RolfuOPT3o=
`protect END_PROTECTED
