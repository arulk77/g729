`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44wp9ApcGclbWBnuIPcYN+HHEdg/BLgbt7PHxcvWF28O
sYRdDugK1mvsun56MF0VLV+LH72/sB1Uahv3sAVkkFXH2HRO8J02Gw+eXGAZJ+Db
UWGLk5/9+8uA35DfCYPkRuF9n2GskL2gJIrpP8JvMtTcGmKnLXJggpVFmuNqPwNI
EvWE2b70gZ88DgChOR+2dBofc5hRhvcHSmQqtFrUX3iLdtEp/CH0PJ5QpTriIzj6
uj72Ls8SHUklHWoHlEOINSKeK/j7ZfQZwUY8gzLoJdfNIhgvp/mqFkUCQegLssbn
yee6jMWbCCZYN7ulAveVlTPf8bcjXFpcOOlNk76WAEEbgMrIah81Zqe7Dkx2VidA
AJG5378iM2Z2UUL/0PgBEOziw50yWCLFrblzXgZOGY+q4XQahqklDG2Ay8AB+CkO
HLSH2krJp76r2C0GE0aGlXkwuMzCeZN4anCDQyx8jmgsjZR8rhR8jnb4CCkjIDQ3
`protect END_PROTECTED
