`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NPqLSXHCclGj04N4flTCnThc6VSb8sit/askAoYvzr8ycn0sFUH68UStwPuHsFZK
SCDgHt5hMMAlQ35UuhbqWdp/vYoe5wW3TIGiyuha9enQv+QG+xst4mOYNyWcg5hj
Ad4nm6Mbbb+q8irt1K1+gquqNm8i9LNqp14Ly0XGHJUx56FQwxPy0gAWivspMlxz
cjmH8wNS7tazfIuxDs3v0E/UPulEaDfv8vnOOcdmk/jM5d7uoCEH+2QZb1bYIJNq
OdSLMYvCzsGlNt/W1v26wJxGp7un06AUSmoaMfzlGmdJeP64zgtofP7XWLstMVMs
NvDDxCMHreX5+ZEGv4zx6Vj9QkNUvlScHK8SrMA7wNc=
`protect END_PROTECTED
