`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7jzQVtGELT+GlljlZihyFO9DOqQd8/h1b06ITFNlCHOq
191M3DsPo0SkRVjDr9zHtwEPby5Ev0hQ7VbYujrW37wNG6vwnHIVg4y1Ys5s9Fdg
/WcPA3pZ5pcJ3lQGFhLcVtOgffcEzlO0+3noKZUvtvlYln9W0EYQ3qrGQRpN56fO
L39XDnnMTes/WBg+qkwioe2Z63Z6YasI4Mfoit2jmpBsTSXHLFauuR/364NPf5j1
YrOlgr/URYs0pixnYLhFbp2R4+98qgyIPF3lcA/F7lgkrnDZ09W4XWF7fQ7a5jqX
VbrxL1Y0jhLSNiSoAPRc97HejPdhcSVQpR55gsieNbLoRz+Rn896ynSkLFi+yS52
G8Z/PiGLwykA2G5afRwHkxNzl9DFpPzW1Y1uMAmoWet/Y+gkg1D2GFWPWqwmNADe
XhKdl6sUdKgCFhPTjpk6JZxOsBwEQHd4WlwUAaq8ILBQXz4koAknOYboGhUaXN7I
0xkKy3iJLXj5J1Nh/Er7/ngj8gaywq11n/EL/p2KdAnhroK40Rif4G8d/N4PHojB
fRO9Llo4my9Z3rzjPIOoR1zobS/SaqoiaaNtYPXdQb40XU5gsi39Iaj0clvj5PvU
LljCFM9b2KctBz5yEB4BdK7esnsXvoZOgCt1Sl1MWIpwAiS18SNCstoKvNz7MbrA
GHXPxdZT/alF6alJgPzoabXvhZ9EFz2uQ54yNn3sLYAaIUSRNpM36fjchS/GayUg
S3FTI6Vb+803MDUVqyYLH3aEOnVq1hejvn+3RJSwV9m6wefgFGlee7bM0+o+Oq5c
WNhqxplQ3WUhIV3IWr163vJhlF1CgFrTp+nj3xwNZWn+vK4xPeecfdCQeKSrAvBQ
ZRm0bgOZ8pPWjcrbABVRPbqcMeUEFcs4RoHsmAX19FqsUJFOfvCagizdFMO2Z2Ja
HUU7O5Q5IubJCvGFbytU/Az8GsCH/lhEFhGa6sc1EAiikXcl7i+Ad7mrPLLa2wDE
V1nP4Vfd3NDE9a8NLgH1INPUgKERWv/0Xvt4qYLd0cJOsmaTE8489h6eEMxjJxuK
Q0X3OiJmzrowmEJ5kfOQ3TW9p7e+uSO+x2HYYsVSRAeTvh7SCu37/KbeSCm1ya1A
NXV1f1QXZXcGUFGVP6lUAbCwiiZz5P0A5gUvvqRBZBE5d3tzno34hfzzksdMfnUj
G/1Lz2Igd5BQNnQWDy4c5Q9EY4397bDSOJU5vLm3fJTKrtaznhAzeTD/eDzKWbyr
G3auSFj6b2AIbe6ON8riSSiwoIlBflREO1GoP79t0a1IsVLpMxpP7iIo+w9UcaKi
58/0kqRBWnYJ+S77sw0yfhpsULCb0hW+MTaJwOQ9qkHjy9HF0toISjg6MbENcLqb
82GqoWunshGR/Kq0oEtg9GYGzPfRy/16QKyRV3nqj5xvC2LlesmEcQbCfNWy20zP
b4Q7x8ngVVVBtDplmIpCkX14pI76y35Qz5HRkFUz/Ef7UEQUwfMXBkLvSlgAhjwv
ALEcAPQl4wMrXKFZmPwAgoE9y46vBb5H+bxZUWHBICb7sDGvJtSA04GiD2Z5KnJZ
y0vnc4NRqtK0g6EQJeTp0DODaW4kf0jd6VGc5YIKKCP+wrGZvFO/sZTkLIdS2Gf2
HlyT07szZUdPAPp3EgWnLFj9XAscfya7unVOPoIZjRjMoK4fBRWWDlkQHayvb+QY
yNkjNlIIt9AOWUrtA+S0nwbQp87gAS52P637af6GbrDwC7wNjZpg1CwxMH9HQc9g
y/s1wsNX7LeeLe9fIkizCuGvNeEuo/nZ0Ag4ZAErCdmsVHosWsddLaVc1KZw2/zp
eY1SBQKdr4Dj0MfDghEPD25OuP6OF8+uD03lHh196GMcxhQB7GcAzsjthQTNkeO5
WI4+GOuaPpla3bvfoUp2Ub68X7ht+IXEu3EefiLkq0tx35qIeFAYzB2prD1r8iW6
2P7jSYv7HAyaLo6/e0JnQFloXvu9fSaViYX9arKkww7wmcZE3Gbe3aV37obRzX/r
o3gM16hd8Ihgy2IobbmPUF7OLgkuh+iPCBlpOk+Dhuxbr95OzZCgXa8SREXbZ+vP
X7AubrEfYuk9q8m2HwUixzaWqlC+5E6nqhM+OitJ6rrYKBxO41PhVOxNyZ2hZT24
gb7dFv/c/fq0095vBvACWwuwLawhnPEL+j9JzQHZAjZV85FKztUqzJgvsJ/xxt/R
nSoAQAPntjWmxivM98sHlUCZnvGj/7MPErNayY6eIoNim73S4D6tU+jqvngkUuqB
A3FbBt8qHCj85uqwc/15u4KJKB7vZTW8f38Tv/bF7i8QU04kHGsb8jmJpzacCDeL
JgG1wC1e7QhUET99tC16V+nh61f9w9FaWauEzLreuMCqUL4VK13U8JAXIFJhegMz
J59SnFkJhYvSV3EJcrIeR4M18Ija+wTUzRxEvt6ZdwCIsPEVxwgZPdZg9tMehM2P
p3Rmab5v6jDn2/oZouVgbdXDmQf6yrlNi1XnjiKGMd6T+zzMEDvIJXXCPNlyd8vk
7zSq/5fxEEx1mRDgTbKf10KcrlnD/a5XQnZMvkvTDwSy6770Yqj32jPjwy9HOnkB
rwZLs1g5SbRSXS1FvLYRZ8pRNai7xEx7Srcq1801nDST9Y0EoblSTmZh2YwCYSd0
GL9LTqnmwo69rnBE9ZF7tdowWndzUfzFrJJLoK+QggjuLlC6eFDTk5Ik2zB5t/5e
nc6kvXQ3Hh3jo9noI1lCzMc+s7MsAGJbg0RafhssXRAEQIb71P1Z2XRYLJRE9h5S
Paa/qwduwaXIh3MCJ5UNGhdF9orPPbvYpw9xaUhMi0wzxomVQUlo7NP9A+Fxi4ju
YbgVURvExlSe6sv0aF4s2/ENafbwiePdPyzrPkb3MoeJo7+pvOi02welnk9Ve/Cd
FcI/AYs2fZs02rSbrQzrBn2+/jy01I6J0fXEC5K4gvoR+CFPIl0p/gY6Ls3CRGXE
SjGYsK29iHKyARGjHvi0fRG9zvmxQV0kyWp+x1G/EGyeTAXQ10adaSF7+rsf/HAG
DgcAfOJacLMEyCm+fhvhC7CacaYcCMxG88fNc6HEjs82Pa9iSA9QZ95jc71F4i3o
afV2smkb09y5+rvTfxclF7NOicy+f18Q5xQTVvk3gKGxnZtAQi9T2UF3VVx+npjC
SbYGiWe7pEd/feBnouZyrDjAn3S/KyQqUBYyyAp1q4Vpta+5/uVbWAFr/bJ9XWc3
VyV4AEUCmzYWCF3PWAZR53CgiC0G8Aj0iX37E4PQ2wc44pYYLojzYN6FAGLHGZ2N
GqG1dD5jBi9mAxjN1B13ey+UIZ8jA7nC3HfhwwW8KH3cLQZdFLGu+Pal8tCNzt31
3YpQvRrBtc5CY2CImm4hQ7GSobAJrIUN7BPpJUogUtSDDNAZyoX8ojTAlCHIAUkK
S2tmQ4+hC86Rzy03NmEMpwcxbXZqXFszYlMTqIgvYBy0TdjQr3vpa3jtpPNa/8xP
Ouaq9drGKeRoYXbzdKUnPoBeSFxmpq8zG8wZ4zPcza5D0SRseH8j3D2aItHOTkUy
Mcz+NwCt9G5ZclTdOeH4q24AP9bgSX9dRx8bC35Rr+H8NhcY3wEdzeBAXZetQcHJ
MQ+06l6PV5+XJIkyqo3KilgvVFPK5NslUNY/uD4wi46quYvunWN9/k9gx050CZbT
m0s5zTCPNg7kfhCSMcnt3wLxsjD0EvvwUPQrux7jAC4IoxEWFw3dN99JO3LHR3Wl
Ge6eO3Blbp8eh3PtsXqXwAY122xzPSBDW3YEVJcDaOHQtk2KEa8Hr33F0M2DeYCB
KMqFXXVCRUJA3zec9WtSHuRC+GHNdtT9/4av2lGeOCYdNo6CEXayXlV5gc3Gmwai
ndNUsFNYx0dpO4CpkcEwcZbEIjXvAf0WHvfyKCpu3Bocwz0s1ZQZ+2bCWcVfFvJY
BKpadu5nn1XVxKkXsXEKHJ888DRLKN02CSnXdM7CBTbbL161XRycEEXXVK5TPkrn
HTi6BTjQ+pvWVW7e0O6BVSp8CAu+wCK76qrBB15LBMHRx/oJECltMe0DRl5jzkrt
Sz+GOWQn0r5jwyGczmliLLlgqiO7ECAPWmZBh1+MvQivB+B4O6XjMK6an1zNCWKl
F1NrNcJcAUeoVD5O+MsU+7v2NzpF4BS3eua0egnfJjE5IvV74HiGPmmrDgz21EeR
O6RZOt+rzumZ6coHoZtzql75fw6+MuGH+WmnmKVGoZ0VAaWrPy2hcMpyUNW3+3ju
w0LAJr9TDpgZ6rexCV3Wcw6jtArxA0wkDBhBU0SNDsd3OzWedL0udxQ1PHvBkdUD
DEgg29Bn+yVARxxJBePovqnX/wnfqFYwm4DC4daoYO5jn8XsZgSZ57o+egv/JRJz
xHhvfkbiwWcDlEEJtpHw4oxepq0iVOMbO3YwbGAngsZlTST1Pq8c/IIpw9onAw2e
uTlr2xRrGC1QyLxSsSfFXmNQ59q2JWQDeTigSQ2LCkKdpWL1lM+tm3BBg0oK00dq
Gb28sEOFsPYKWhvoqXtsx4CsmvQz5f41KwV5CCKh7qq++cU8mH+7qgLxR6DMKjzv
by7FK1lo2QEhZn4lUXMPUDjxhZq65dnI8EDDSk0jvUSxyKWT5MEizMzElF3m5HNU
MyQhcv7rBrATop2o955Ul44vhG3aUTZUmXkD7ryLXSWmVqSLHyk0X+7C4JVaBn1B
xQkudhNp0jhKzGS44JhgAhP7/Gj+cpLRsUJQ98dCRj+P+4bsE39Txt9lMuFwGvjb
mvPkXb7NnUBlozx5IVtZx229N++qY8YspODGFh/BnIGLPrAH30X/YPKwWxY18Nb2
wKyqDKN42gnxCwVXEZPzjf+iM4xv+PjRyXxw6fTRfUqP8u8HP9E89BPQhlog5lvR
cQ+CG7sYhYEd5bKaf1jXZPpRPS7j/RZNQWzIt2dbeQxGoWphSkMOvC9OihP+o9Bj
fx73iYhI2SC+t1L3yNqn852RbqmK5mp/B1hjcyOlI5EzeR/V3NedF2xcZBXlgFX9
l7vK+AfNx+kLZeR4VJ0hSdKtyzNWocXQTscVTOCFsbrBZWpctvaGaMrHwcEOS2Ov
NrirfkDXMdNOO0tS3cm8IrLFsFmZLKmhgsE3+4+9UD1CTA+jhmBe26OM0MO0IKL7
5e3j4Kdzt03/zGbOeufmn6zKpA7Tw8IBh3SCoWB322noibncFgjP/GCmAghzvU9x
oHOVQDe3S304kBUwcl1X7h/rSeMKuK3xwXacUpJaIkkqBK3ETUR7Bk1tCxdeB4N8
WDupliJkFpqY+am/DHsAOQ6kJ5dnRui6/nc89vRvl78H4q0lQCokQ8vpDutGr+Ol
ct5XyBGyG8Y/7nmH1EUHJsiMi/FkCUqgzz8M7USvldKVcMWC8rygpnSFOp7o8R0H
gwHdfBT81/XpKrVNL+R3UFhWv2izYTQVcn1inxHxieWreF5MQNa2cS0+2Lk2jQqB
MeIZZhMowICVNsb9t174YpIkUpu+MM4YhojPorpEQFTbviOX6csY3dkCYRcz9///
TcPojORHNF3lIi6vEMNyYf0Gm8g+vhuLFdUbs3Ldu94tyXZGqIzu46p1VAwvE5Tv
p8IeEZedgFIgf3xx9urL4lpmts82aQCCI0EGFUlBidFZen+RcYO0+M4dJepqvmAj
OON/4uxneoczmozkurXh2ycT7qwmTjDBxAEHPQpz0QeZOQZTFSMZB3tLRYy4EUqD
Wzqsm0hNyS0VpZW715NKxkAck3jhDqb6Vo3SS8X/2wvfjTseYFvIc9EjjczgUFQo
X3iytywKmNhwjTD/0eGd5iPqvH43k7bP4m+AoYPMFHmNKYVQMa7QaxbRnCPFftvB
BxjQVYvSm0b9wKhrmxwosStyS1yLgXK7tx53M4yrqbWLXOLNZqUB+Dhe1nrXONLm
6JpzIPAWx/pSSbyEYHM4OAwUfS/jzCqsDSGMifEDLfBOoZ0SPWDl3zrC6FDnW5Qp
uYJ+SklGbalm38NExqP3G5oXNXL1aLloAbJvmje64JYVzdmMf3lwHaCyXF0pQASf
ahkgu5hH29PbX8mQE79Bsr44LRaKHSh4xtmPKf8iiqB31NtDMjVwC+dykBEcRuOj
Xzt6o+mM0NImkw9Z5E44tUbxANiSw5+zYuQd517V9LqcFwWW7ctZIoqr7LdGclec
mhtyQONce1rKoCvZaY6a597uKEyrJk/pgcwTwg7DabhB6fLEH85T7TBWFOJfNAwI
/G8nNj4uy7UJNyjN8iAWN6JgLAiAXAoLocqsWdhd1mMOfPsMA21ok0y5BOF93Qmj
Bt7o88xVr0q4nF6m9swUbhnVIolVADFfMi0ldCTZ1PdvWUtwuXBkMffsPubH2rgI
xynTRxQwUCw7BAFTqTzB/sEyWOFmvYqx64woF8J6TfT4ufP6yqeRqmT++as405wr
QyIwYVdPKQd43jcpwXV8CHHMa+A+N5ip1Szgv7ODRqwwR3KgLzvdeqwBqK3mbHw8
OAeFOjyyOW5tZ070tL6727I8TfK5dFuTVLY8Xhtc4mZdJZYzHuBNnI1LcmbCoXra
BRdZ0Pts0o/X5ZJRPcGYflTinFuhGPNMO+Fa4ClsDrt0SgY2FNtJkv75VeA6bYiQ
RLPPck6XMQVycWGSWzNXFy2Q4gHYwlxTxwSyOiU9TcHJaEr9gNIPT+aaR5NKTjTT
xS8ldNt8KIOmoKklQW9SgjzPMMXjA1WeuR6LD1UtHU0KjeYxzHTRC2whW+eafTpG
ZsuKPDZdIROQvitjQfozDcmSA9yzHY/wdACA6a7FU4YdfWt4+x/v+V1kYPP98ppc
vimzV3O5bDQtEVXyGGQO7ysFad4IoP8S468k76jW2LtzkAxveT6y9OSc2qTUuq1z
HST8HV2bQjGkFgJXzyKLFxIr0MOR5Zgo29by6RBsCyRWaiJkDDeuYCvarsF5usar
Wm6oD6Qe0qpw9x3dOGfWjYX6V9fNcesNU1zeMffqb2Ua0xprkGrpSsfEWQvYzf4x
S1qIaI0KCYjbvdoIHCRD17zP+NbAYYgQUpko3ifEIAYZMmron0aere0MMDPZ8zQ6
fo9GFoGzVqcECvJKYloDH4AC7HvhIXQcjWKUnHATr1PJ753MgKEfeY+bbcAen3Vr
nSHkj5aNSLR4gOB/BYe5bF47AxIpp1ZHgE846RS3Ft+ICKtQpjHGfyKLMa6LpxUj
Deuc+79Mn85XAEtqip1JsKy/HGzo+XjxIJnmTrQMjfy78gI9pOPOUduhVkdib+N/
RFc3OzUPnC1ki/HTaRc1pgiNoXABL0JNyBCRgo5aDUrjYniSK9ZX3qFqPZHq4sW2
yUxlNFtQcy1dz+SmlV9WBeZT6xpVrT40SK71XCS7et8kIFGLgLfF6lnNlDJseCrb
qhgcnpcspRL5fZM/yMPDDIXK6/Rd+r3JponQH4QyHxlHRxETwuJMIReT+Xaf9lQH
00OIVzIvAmduFgEKABqRn/6459Zs+piFskFlAqXAHhYh5Rbo3/krQ4b+wbZLEnRs
z6QlxTHALmu6Nqyu57Ww7Ia9zL0vd4B59reCjhrcZhm8TVszB+KMPix9JplXsdF/
moTXaUSvu6JFgFWQgXLjzmUn9Jw80kB68LwtiPN8Y5qeFhuyYaoxFbpOnkhRu1Vl
vwK3cgxXn9jjPFHCHGwFZ9a1y+KWY1UaLbjoOTyESbWMpGGy/JaGdN6oByX948y4
KDdn0zQExgjnZGvUuyFh9FT5Bb3p29n/erL+hADI+8iegKPNT2symIJREgzJHVbt
Y6SouGAI5aLMKY/IVY19++Afsupz/w9ilsh/xjLah9rU64qkWeUZq6b9WLxBr3Qs
2py7c89ch6j674lDWpsfLtuzxDvkZ7xC6zBaPnZ/X6xPHF9K9hONk+oge1N09X34
Agm5DuqK2ePZjCdXQbUGQMqDc0vhHwXIjia2RqUMdVREL3oCZbjNER1lOpge7HpM
f9laAgCnQG/PLC3dLALuhRpCXzAXnNKvKnj67yiC93SlouwzhiBaxMXLyFNZIDDR
oB7uKh0DrljCqiKmLBoaHMCKUoOhjRD20f3FhCnSVhsosMSgglgZX+zflpWGu9tw
68QkPpgRjGh5Qh1ZjJqT5ij33eZcYKDBysApYtczmVnRSKq2vnFOIs82Pb92yfrz
zeG/X0F6g7p7vph9Bum6cQris/mmekQITjEpjPuQqxgbiLT736q0sO//4w+EWjjX
RnsiyQPmrN7GI/KPYxzy1y+XHPyWtM3eKJeBIpkFS82sAk6hmGm2b5pHSgaHpG1Y
F8UDt+4wNQT8bz6f3K/8kxJXZd8dtXAnJgZ0AY1mGO2JGTmqUbUl3eB5Q62f2FAm
JmfW3HIYqCHdkQB22nDVNNGFZC01qXohvPm0ZSTNP6dKmBpaC3vCPQxTINdM4h15
9RfgTUCnVd1BdAiiWpEeR1FgI/fNlYujjc4qbCU46LQQLkWSN8SjOsCTLkfClUjE
4OP+gM5y/BEBTDPEKykq54uEQJ3p6oWlLPTzAlIziyggKIDukk4+dN5/b5CYXC10
n0uW7Foiz7OD1PzP9eRXgen+Sp3347F0CUzOt+i24omrR1OpMhc/Iv1qJCs9kKbv
rWvCbf8tpyxx2n02aTPI1YNtNW97z8bZ29PrrqLCKFSXNfzSR9Y4qJWrtbmKGi7w
AEjh6eDvRqpvWmyJAgGAcPltWsX+Y74lyHv7t9u8SB41E0e/SdxQS6PX/XcoF+2p
+sjGbxhXcc4ADwGlyXwz0nAFnTpzGnSjoEaU4Qa1jJ4qlBGyfY8NOScRUjj1pY+T
Z5tUbwAQYl3n2FRTzej/j/ranewy2sk6F3pUSc/HecRn0hzy/Xrh229Zuc4qnMrl
ACqAbuzVzTfEDfzIudKgqXMBKcnpi95b1ssVAkjseP7NyfYvWvafxVP2foZ5c6Xj
17Rfzggv2OMZthroMCFODgx1IVjR7E6hIb4G/ZV35jW2iU/wd3f3ig6dXMQKklY9
umMglrXuhkECeQiZhbQS7wHL6KwpFGQFLHH8CH6mG0617A3erp1qrhPB32ES72MC
g77sMtmV4k6ObsPrTrj7dp8jQbuKuEcErqOw+cg3wOjF+E8Qmb/gUShlUaQzuQ/u
Dw+vCxNUBHO/QuYp32Gh07nn9VUXP48Nq0ClxMaPAH2UGkfa7AQsG6eVhzDh061o
Vn947dQysYMjS/6g6wwF+Jp5o0cSQlQ6XORaeKpaIRFi1rukty0DABqNUiCwGode
Su51xHRXoL/2cr6d3OiePqhvWh3VIZKvRSNOParuBSC4+9KLFwfrA6220KIXLic9
1tlGlNbQqO6T7q3r0SdYW027pg7AjZpUZMAYbY44cNGT1pVqf+DgaVqZbYhiw1ay
EUAvl4Sgj+cqWZKvemih205hZHXGfW3UBW+zdKcho3z5u3yqB/ddpu02VdWLsmNH
Rj0IlWKm+LJeugCbv2+fbqJ9I4ryQCR+ccjJz6l3DNtvCHx3i6kfcSzINdWuqFdG
r+tyWI4FZ1hIpBkBKQ4haA7S02ea48cRmg85epKV1KNrgiyeUShnBJa3yfGdE+GP
j0sI0fA7VRya78qSjZ+MRSlkJJu8DrEER8QGkoDLhIr5z2MUS9EpsYY+b2gVRj0e
5d3mzGLAxOqDkBs0rkkY1sBKfSMRRQd55h4Gh+3pVFNQC0VqbrbpsKVICqlWU6xn
dSOzbaFEx9PRai4s7JR0f4UWgJMq8qzki91VqT2VZVqUcHBA5ydFx2uGRCkcqDhj
739HmUqbTezUHXPHAngKjq7wfvToWicDLPEFJeMJv8M37nmZKbz7jUHjxpzz/ivq
oncTTz4+rmNiHqD4w5D5L2+ovY7InN1rHoOhklDug01vBlXv8G52Gvl/GtnomY4T
886C9UOdTeaPGqZh6lqN4SNZlLs06iH5g5AxpBKS6TC/w3WhyDmPQi6Mq2/PyuSZ
kP4MDuBMdDyd3n41VXPP3PgA801fGjhDmqct0MiXc0CbSdgmMJNM8UTIUwXkhY3u
SfzjBRgVhMQLueOHhvxlXP7FDfPm8LsXoYQ15mvUcuuWSPBOpvhWV25Oq/yGbA5N
PQTsT3/q2yeGTzfpQFICV+icBja7i3KtpbK0b4/E1TfF3SWdVuGqMIcIe3HMuNaQ
rsalO8uuyklEkWSXse6atgvrfKGQnC7g8GU0WtbsgyH1wDRCzJ/M/O4nDEcgWRV0
CPbmCdRgo9ghVVpTOLyaz41N8rka1PGFZZ4Ew9tNEvHKhEEjg/XbkkjnQlO2VJuF
SEUcuoBOJzslsLnqJF06sVndVCliXhCNkRqrCdlufLH7c0/kc7ib2uLNp/fKAXAt
u8HkY1StF04y/Sq+xdpd6icL2ysA5xk27mfre07qKqkPpe0iXdHvIcsLoTFzYIF0
UKdjY3J/UJrpnkXTvI2CZ+alhqWlFuX+TVHkJYfHEUQTG9BlA0dA/olx++IjGriP
qwywzo+B+zrCg+lXwrqsm0/Nvez3XjAxAYeCQQLZopJmJ5u2pxHJqYf/3MhN1tHh
9O6HbVSolVvXUtXSLGDzYyIjG7LTUlbSeWZH41YrRYg6iX81Dm5CrIVUSBjUPAi3
iLFD8O38zFJSblrnp00J24E0Gb+H+ruFlzb5gSofL5T3KyJ4EoeXVL/sFkdbjlM6
6w6bPL1y0JX7I4ExeAcPHioo7zVLjm1vmRyzWUdsHnhZNO0N0nqefFHaJaq3yy1f
hfQBKtRKc9wFbE8wtqGEBgLW/HGjF5MyxPZllze/z8OOVxeZOl9ydP0x9rb0MxPC
ATI4dvY8iZFRT0n7v+gEsvDy4C8YE8/FUpwTRz7L3fSnS5UeGFmaITa4n2V+van9
6LCM83ab9HScJ+drkemzclwd5Z5yJa3bpzsx36Yh7w+hcGLTLxD4IgP4XZcsdCwZ
Ms0cmgNZlMsplbYOq6nlyyNyoGhr6iOUcrv2i526CIqJRRIKbcj1ARKg8KtMDlh2
BilZH7iKlJb02nYTZoFM8mOVv6E0hMmhuRiW2ZUSSMD7ug9p9aYKzZHt6FaKA3cS
2eahaBxf1IAwhlPut5EtZxP65zOIFmYDxFYlLKrkSZ6Q2ubpMbvrOHJv5cfOD0KK
awSj1wLDNOR5IocNyqY6ZYhZFGZXdvMgnDGec+fHkUyOxTDG0FjIjFLG2MIJwFoH
52HKoIc2A1yuCqC4FKo2A0I5v6LMC4RXNHzmEvH3k+hElo+VmHU/RMhPBwUhftMg
MOVw09Q1iLsHEgXx1WiWuEZm5AkkpJY2T111f247nKvojaRRhTn6H/EuP5n0/0qF
6O1TuAkI3K+QsrR4i5qBIZ5d8GLUIrq+wxaKrGGiPrCvZPO4dw4areRyauSZf1He
TgXduemT/wX3kbLHDsVCmqpCJx9NH1EYq9QbcMOSd8JLpN88o9bMEo2omQJWx8L3
m5tSlj2bOzLvBes8vN0jqaH/wBypX3LzwCp5/med0RVKsINUjVTtrcHCO3DyOSJj
Ys0oMCtN/eSFFmaLyZ/V8ZbyxEiIHkWDN36tg1kxCpFe9rBiwhGYIste21rwLeQr
3z3s7dfznC06OvAk2yjwNA==
`protect END_PROTECTED
