`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCv2kJKYfn2LaJgq2h4cxTxPnxSFaZHnTgI372RyFHAm
+N92HgDKFVWVXzNwOpA5twgX64Dm8S/c5V152qYmnk5kzYxKfGeNwK7QNbFrdeIx
Z30BQSjbxZoa7aCPSSVoyhGuP0i8mz5G8/D6/x4aKiAqedvHKbKaBZ+b1H2hBMoB
p/GQ9tIV+U3jhCemU5EkbD9sKI0AGriP5ZnkQPLyj3OM/MuHUIKGv7rqTyPxys3B
P7P+FEW/Oie4Ho8rQw/B7jI7qGkV3BQ4Rn6LCkNHwI0xfpOT+ZbkfnfDbSpgYODT
Qk9vrLjUt+Ui9c+lw80cD5tO2DqSytNX3VS7nOz2ElXWe0egBO9pWaka4UzdgwrW
Jc1EXN1LDGu59FRPHjTqgXGn445rN3GBL38OmvyN0T3yXsEwswUoJDXn6cMB49as
da31htEvQSVt5JNyXS4VZCAhFhUb78jQEBrmKshZqvUx4M2AMiM1c79mzga5K4LA
Fuz5FfSbCGhxTjBFwDXcP5BXUzU5N+hUSQcR97XX4seru4kq3rvXl3s/lxxkszfr
j6ZEoXRRCxDiel3mrZfxsVIhqW8HGlZ83ev3YLk7IGSJ5PIoVG1ZkXtC6z/ZE/bm
gsBqDSpsZCkrfc1zmMn2vDiGMXU6CKh8+FphTevjFa9PFGUyP1YT5+cCuM85WU+y
NDvETA2gJruM9jBgCPd1U+Xuu8ANsw2bPx1delPW1XD436BmfxYq8Yea0MLPDt3c
Uvp/LJEovUHmm05dbPTWzZcdS5e+YTZ4pU/cYxYYl7fzegKs+gtvHYhMIUi6/wPX
llsii6Omq2hga4hAsmtqH+x84USWbGCIJBt3RClpNXr0Ttvt5/6003twiRrNkkUR
lpYsBQiutkfbx/2imeFwNKXWg0y/nv6sT3Bz3pWHb6ai5svcmYquzABJIZC/UHo/
dH6dOLTT7Pqfvyj+zlkSFTb/uBeZZKSEcvF8YIrTXdH7N/pCZsG/TcE5M3by0y7k
PLy+uH8ZKoEjk3kO0calNS2PQysAM1PgfiiNEQeZbspgTP017Y1oUR2XEWQnALUk
5D7QH5TMsL25lVxxStF0g/akkJ4C+5dOK/uzpayTtaFGSVrDE8QoaPa0p2PYfA7k
qBc9SzXDkeiNEvzdxmFkcbV8BWQlX1/ZcWQ29mHJ4pU=
`protect END_PROTECTED
