`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAZvv2/1QETxSi8/6YgPEMoaSaboq/FcEDuxD2rLSj6Lr
fqCrFOmIK5bRONi7i35ltH7mUs8Xm4m/+8Js+1w+f6Oi34yJgWyiV9Q5frNoTpBy
JUofP6UUu/f5FpC4EEVF9TwVFIwxkwk+FyM+4nYQDlNf+BvbJZZal1KBFRhrgalN
tycGLKo79DZbZ4fwO4EEPMlAS3ClkE27Dk2U6XxjhVYUWOAGeDVBRDi/3r0/F6G7
meMcWYMg0dt1cTXHSgMZlfVPpVX4+JSMwtzVFCofnYshrrYyT5LNSy3zWyc5Megk
FSNe/uwB6Yisf+6/osLD7rsO4QKs71bgu3MOl9Z8CINmFiVST2zp/2nsfwRweU+8
k99jw3ULEjkXyDn81jqfTLNNJnezUQ8DKBVF3V7w38j2p8jw2NQNXwqSE9G4Odr8
oO+8UGeHhMK6toO8fh79ghOEryc7tffYEy9Nak/16TQhPiiL2BD44Q05MA49lI8Z
HXuBXnTfxd3IzRBjIGZR1wPW2gQESITIokic4xKYAOmZa9CsjvGKt+AZTnjr2V9T
beTfaTHd91kyeY6j64NSbeNQa8/aiWCGlSgn2o7Mj4MhAiq/1+2KHs7c5Yk/i+Yf
nXRN+j0kriUyNu7CUJJ/zrTIJvxqiwmrdEMQhLTvp3Sp5BAriHff2GoJJOa9AN24
VZhI0r4Mg+4DsyhmBHl2AE5CFluWKv3MphZKhPCEPcgqE7SiZdci8ljI6Oo7vTd3
fbZG1Ua3gqFc/ZBWSpXYPshifMqAEs2b8tdKtYYCCbpI1SGAHRDdtAd9Zl5l1lmM
vjpnRWnXKIbsmn0cYkUaZ39LsQrgai9k5dhutCcgXG69Oz+AjQJS+PE9omcsLckD
k/McBPRBo+f2Y7IJsCeU7D9+rlvUhNWItVKLAp39e+h0VpZk0bUIDCPIm8RqjUat
p2BGtDdR6BKP8EKGRUCzZotQ/xOMahnOkfYhgg9heyKXiJFsS03b9axP/AK3y6lc
s3cjSk3Hh4C6PS3t+I6LFmcksW68+UR7JpASRnJhMDeN91GXwznqiHQAwpMYg7CZ
VCMn9hVIqD5elJ5QutHyoRWGUepJ0DZ1rpR+B/BCE6xV3hsJ/21t9JJPLmaryQJm
40LBU4V4kLsSD/2xYAgzHYRiXLy9awoS1k0IJD5FTPxmBqaea+TqMq75ujl4r1G+
35IhgcBvSK10UL2c6sBHhN/iyoVBmu7JwxVpOlfJR8LL/aVB3rCkmDyx8Qb8Ei3y
jqdOgSp6XBwI2LsO4KD5ahMtAj5SztuJV6NrK35e/hxCH8U7FEkPrQ3AOf86q9EE
F4dBQlrwNAdPzq8UN2elDrJPP1WxrMHc/0SKiw+mtw6FO3z4TU8kaVtWcQ7iN4+w
78GpdOOrI7Sx+PAxkQT82g==
`protect END_PROTECTED
