`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH/O+tLJjszsdX5aWU28pYLiUhhUOfRJgjBi8Cf4OGE4
mfZDLelgH/RcgjmAtr3P4vuQ9LFGNWMFy2G731mcFfyBX8CIxT1EtDTAwHb6QJRZ
0mb7y/7lSLjvUZjLyMG8v4ABpgrjKd/BqrdnVojamweth80NqOlVRALj6a2BOxyk
R/kODosSyMzCMHbu1EINVX8audzs6IVO4TmaqHhzWzWxHWqZPKVNi0FruEjW55+P
H9ZQXvMplqcKrx7ntjpY0GHtslMH27zUYXFVum+NYjElKCDyh/uMJ20zBRLTJib6
DWGoPXdMZiISyfX+wASquNH4mlJuQoM9Nv7MMYPS2D/nllnwYzWkyjL6lwvbQlq6
d/L6bW9tJ0gM7nCnuJwovxfHvisBqyqADSyet+qHyiKvCkOSJl0quMu4TwJityfY
Xro62FXi7BFeWRCxlzC3hL9h1kjNjDAekNR1G3r7Ve+lAA1pdb9tCf+DGDafcPUx
c1eJ2e/xWjnmEnxtbDhJmVXYIxIfJKOHL4ma+XPUo/x4R8ocVFrnBunBqNGh17hU
hXFwJ7sgDCZIfyY8vQSPX+UiXJxdlCGayAKJoaLJtNIPE71iX/ImSs50uJIIcEHl
nh5zqJR8VYH7uxhbxywVjbCI1ED7Q0hLOw/zFipYnRnt5Mrd3sj54qI23VJ04PvZ
PDX7BniSH2pDtmTIcSTPJaCnCDe3z9rgOcJxTD4/0tBDuXbfUlEDu4ajf6uX32rw
4+/ILHL6bXQ2E8wxRZZhFzeEPrrMITBv57JlYtKLIf6zkOIpVN9b4BI6ljjjFx6N
sgXAIDF3o/pAi9XzwomcRUBixPC7V5Jrtvz4uKoGaHfJtL/oyvWBqwVg6my0oBnK
QP6qVvUU9gvsPVCRlHoPZqYvNZuZzL8rwFCS8PykErByyvTQbBZJt8HPx9MoOBo9
IwAu9q5MDD5+thU91TjwbgEhN73KZ4R2rQbH3Tn05eVdyvWGabyjNnnA6A+5p/gI
aiS7Rky6Whu9JAr9QAGzKnNwkMO3U1flZpGoNP8xoEmpVB9stoIzUwIGU6f6KIDP
/UNm1qqGwzzw9uGnqW5lopC75++bXPwZ1ldvl1TlQd/g8pzda02/cr4b7tXUuUPn
lVEsMVOzi8sxr9fKXLItiX1F6I3sJ7iwyvK8wm3opKrHUabqulu1gJnZ8/taBb8q
i+WtWX3zx2EY+SYbCXUVlnQCPnUvXm+bYmhLDVzqesAUrj3+ycmoisPMkbnOtCAn
jm3hxybAL8hI7uV5ch3qMNfUcJbyFtoeRXFkwZeK7chdWjS2Reve8mDne1DUrMV2
4xox/XsrRr2aW5wahzjUjQi59EyMqDF5CGoNzaqYK9hakbMCQYEXz1Ehn5iHKpWt
J73A8Cvn289Xxq5xHRKJ4kgUnQEHMtMgwA4R0ZuqAL4ArqSbO+uWgmli+2QVX1vu
yai5qrXc4WkIkOXvevQac9L0tKbRSBs3tym4z8mZAZGfJ7fvJB5g8QjSKPQcZyDO
OjOYOjOrRnvl2sVAZwpF9su3TTaMjDC4o4SUbrrGUS8LZ5zfiIK8sxMOSeSdhcAJ
npyTIy8Zml2exyFwTuTqBqFXal7xvX5u2usquBPgPRzoBJgIVHPcp0TWZqxg5IjN
YncXaVJMvfr63f1J6yHdvQ==
`protect END_PROTECTED
