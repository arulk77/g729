`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MA+owael/g72V+l+ftZ9nDWfKd1j3n3c3BIGQsSYWi5vp6B7Ph7rV2n1Lv4R6ZD9
uLJ8rCHhbJUWkkXUqBVvz1sBRC4XDHC7erBKKFJ+0ZzWyX3zxJIxfmLp4vCGarsW
ARzJo94RCcfDoDBImNgVIZUF+QIIzkprJzfxcNmOcg6MDxXb56q7ogxcFe2gnwMw
XJjP1YOAyzNIj0Gu9vnGCRQ2lnct668nKvqfOR3S/6pB5bMWEEhEHGEo7WKPzT8/
ep+y4erIXskOkWB27uqwPED+1lrmrloYKILpizSaGmuWq9kM/a85ycJJUq1W66Nf
`protect END_PROTECTED
