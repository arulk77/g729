`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wjyJUspfl8wHnBau9S792/39JGVddvHVimbP5izCIcC
mfW9hBEignEKOZKO20hsu+QY3MDOcIH7VMTO8wnt/4xpcxyzARjK0oGSBJ+Uy17I
oU65COMqO5vYdyvnNB+9AQq5+/Pga66aANNaTyyapMHtOEXIbrdI3A+pUC2A4m/G
jWtaERbmoWFSv7spSHi8/HM+WRd6Z9Unm0tPlESwyqT5jYayG1oplDXngXYNed8W
HAbK7QdgdMq9k5k7vbsxNogCT5Xz8+WgG7OEGVXbbUccpFLim1B5LARmqDvD7srr
MEngIADD2iFsF/TxnesiDDsr9ByNnkniOy2K9J7cxUy4xof0P4bVjudrDG6WpMVO
SiM9gQqE8mzRAWGNoSQq0w==
`protect END_PROTECTED
