library verilog;
use verilog.vl_types.all;
entity MMCME2_ADV is
    generic(
        BANDWIDTH       : string  := "OPTIMIZED";
        CLKFBOUT_USE_FINE_PS: string  := "FALSE";
        CLKOUT0_USE_FINE_PS: string  := "FALSE";
        CLKOUT1_USE_FINE_PS: string  := "FALSE";
        CLKOUT2_USE_FINE_PS: string  := "FALSE";
        CLKOUT3_USE_FINE_PS: string  := "FALSE";
        CLKOUT4_CASCADE : string  := "FALSE";
        CLKOUT4_USE_FINE_PS: string  := "FALSE";
        CLKOUT5_USE_FINE_PS: string  := "FALSE";
        CLKOUT6_USE_FINE_PS: string  := "FALSE";
        COMPENSATION    : string  := "ZHOLD";
        STARTUP_WAIT    : string  := "FALSE";
        CLKOUT1_DIVIDE  : integer := 1;
        CLKOUT2_DIVIDE  : integer := 1;
        CLKOUT3_DIVIDE  : integer := 1;
        CLKOUT4_DIVIDE  : integer := 1;
        CLKOUT5_DIVIDE  : integer := 1;
        CLKOUT6_DIVIDE  : integer := 1;
        DIVCLK_DIVIDE   : integer := 1;
        CLKFBOUT_MULT_F : real    := 5.000000;
        CLKFBOUT_PHASE  : real    := 0.000000;
        CLKIN1_PERIOD   : real    := 0.000000;
        CLKIN2_PERIOD   : real    := 0.000000;
        CLKOUT0_DIVIDE_F: real    := 1.000000;
        CLKOUT0_DUTY_CYCLE: real    := 0.500000;
        CLKOUT0_PHASE   : real    := 0.000000;
        CLKOUT1_DUTY_CYCLE: real    := 0.500000;
        CLKOUT1_PHASE   : real    := 0.000000;
        CLKOUT2_DUTY_CYCLE: real    := 0.500000;
        CLKOUT2_PHASE   : real    := 0.000000;
        CLKOUT3_DUTY_CYCLE: real    := 0.500000;
        CLKOUT3_PHASE   : real    := 0.000000;
        CLKOUT4_DUTY_CYCLE: real    := 0.500000;
        CLKOUT4_PHASE   : real    := 0.000000;
        CLKOUT5_DUTY_CYCLE: real    := 0.500000;
        CLKOUT5_PHASE   : real    := 0.000000;
        CLKOUT6_DUTY_CYCLE: real    := 0.500000;
        CLKOUT6_PHASE   : real    := 0.000000;
        REF_JITTER1     : real    := 0.010000;
        REF_JITTER2     : real    := 0.010000;
        SS_EN           : string  := "FALSE";
        SS_MODE         : string  := "CENTER_HIGH";
        SS_MOD_PERIOD   : integer := 10000
    );
    port(
        CLKFBOUT        : out    vl_logic;
        CLKFBOUTB       : out    vl_logic;
        CLKFBSTOPPED    : out    vl_logic;
        CLKINSTOPPED    : out    vl_logic;
        CLKOUT0         : out    vl_logic;
        CLKOUT0B        : out    vl_logic;
        CLKOUT1         : out    vl_logic;
        CLKOUT1B        : out    vl_logic;
        CLKOUT2         : out    vl_logic;
        CLKOUT2B        : out    vl_logic;
        CLKOUT3         : out    vl_logic;
        CLKOUT3B        : out    vl_logic;
        CLKOUT4         : out    vl_logic;
        CLKOUT5         : out    vl_logic;
        CLKOUT6         : out    vl_logic;
        DO              : out    vl_logic_vector(15 downto 0);
        DRDY            : out    vl_logic;
        LOCKED          : out    vl_logic;
        PSDONE          : out    vl_logic;
        CLKFBIN         : in     vl_logic;
        CLKIN1          : in     vl_logic;
        CLKIN2          : in     vl_logic;
        CLKINSEL        : in     vl_logic;
        DADDR           : in     vl_logic_vector(6 downto 0);
        DCLK            : in     vl_logic;
        DEN             : in     vl_logic;
        DI              : in     vl_logic_vector(15 downto 0);
        DWE             : in     vl_logic;
        PSCLK           : in     vl_logic;
        PSEN            : in     vl_logic;
        PSINCDEC        : in     vl_logic;
        PWRDWN          : in     vl_logic;
        RST             : in     vl_logic
    );
end MMCME2_ADV;
