`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL83f143TznEJjAt1vHIvZrYQZyI3sM28y5vh3u/xU4axk
BCyhUPGWGNw9mQ3Zilohwe5f2C1EYHtwScQmPecdLkjn97pY27g6u96IzqKlUH1z
4eButincYc2h5pTapxDvwvX5MVVEoOEPfajYdG7G1sFQviXU2tjXsLuLr1n9v2C6
k57lxU/FlbfPBW8Hanle7B1DGNLkMsDZY8ElKebPBUawLgnAySndJoy9En5VB3Gc
AZnnR/mRbGJpH4iTif5cJ9apDx4IFmsYsKEDH324TnlL8TiI1CTFGwMdf/vgyIky
u/V3Ym2+EA1RRQcO3pjnWs/ppWSdty/QZ0WIt1Fpef7Q6S4gXdMaNbDavKiM4vLe
aipwC6j9cKCwe3OvDHr3V586vd0J+RXKkHawKDGGgh23KMIPbFE1ejr2VEQg1f86
xcJWg7DMJXgnQP2As83k4ggLUpPGJiVFywI91tst70jMhbMRyOW/q+KDFm0ev5wk
nb7ii9VUPb/WIn90GcsSK/uLR3rTV4N8FBdM7Bcf+BByGqubgFJe+k80T84O90RZ
51kQgwefIsVQCZQqFE1TtxAoXt2E4BJz+oeaRsRQWCu4ZwlINRtVJDHaKPu7gsKY
Uo5uS3ertxLtfVvjZG/bagtrRI/df7fKj6pq8yvG7qBZ+h5nwc2mOETypdTGfGcI
oR24Se3Gd74OKxs7TQND/LssnTETiwYJMyHUsOvT7WSMnb/b6TSSgIJCwHtk4IhZ
8V0lkW30FoudAskeX1mvEqvz9u9ETkOVQsu/fE/sBFGxcGf9hWJBULiiWUuH9HUB
qYNpDKU5xmG2bexghpUwdjEbNx55nhztQOXQWhB7sikjewoJfzPldukBLSrlavgj
+EJui0Sg1oDp/B924FPpCI+gdniDuQPiysDv/olRTye/XGyhyTrQwR/G2thW8omp
`protect END_PROTECTED
