`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
yewlyEpVIiyd4+/50YMeHaoKUPZyaF2rpkhAJC+ZKj5fofAvf5tsCI7DaTmSjzgi
A+rUNuY7B/vRF8sxF7X2lj7dHcCSntL6mJRITqC7Zrnndc+NJyXd4u3Q5aZARWOn
rG1Yh/PHdFK/0JrwXqCEepFqE8XMts7t5nlt9zX7DSx7HJGxuD11fEFzthbrRM5P
tC3Or5x+Wk8FNMGH800IIp/P3MziRxpKO3Ic1QfjHDKXESfrODZdrzBC5MyvVlLQ
0bWhBK8UAah6Ve1WpYtqbeqhhdhnut041kH7pAeDRbHImlHp1Ci4/f2oJ2rZD3KJ
PEL3oI2RpoSIfzaB98Lie8Rp5VXIYNetViV2pkzlM5ppN/X9tPHNAaqCWpTSeRIs
VTIgINYYA+sh1tBs+biE6aY/kGcSoFYyMYDbx2x4z+sdQGusuZhjq6BPHNYey+BJ
gcMwouAr8HtQF2QB/cbke9JBGAHYRAW1m9jSy+XLGuiWVaxZkuinbfJCjsAzlVAW
xEV0rdxhUEYjCQXEkYhkOpdIA1ak5BOPJM6n9QJ59Y0dmi88BbB41AYByMjkz6My
pbEQ0dQc4SgBKY0BCTpSl33L9ALzxwtR34fHNPVWU9rV2x2fYr3PRDw9Uur0cnce
gd+uQmYw+dwmEOlXOG2/1/vQBL58py4UDgCZEQcgQf6WkwmLdMeEql+YXwwecZlJ
3DHJoFLFxWJDki37JFHbvJ4Z73YEx3MrgEonaRo+0Ujwjj3mh2BhySzkTGPMUKZn
encJx9r1vQdEdUwfMTWRBvVT92jdFWDzWvDXCkiHtUk=
`protect END_PROTECTED
