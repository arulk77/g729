`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu482yvo+NxSMwifwOIfCSxPnOPmypFztLLj021V95Lqku
tFTO2R0kEDgcyi7iCoZNzBLnFAbP/uh09lroJC5VieB7Uzq1T6wifOjFcSWAJnll
cKV/FlOiyiykBnjpE48KrfSWuXXDq6hAtf2ppk9IS62ZPau9GxyjQbShS2sVqh30
3HbEJz0RTQwGS+pC2JUNPtLWdch6kbFoLc/+PiribMu1hzSOZat7EJRtmSNq+7HO
QrxGAgcIkL1d+/xSJbujhk9gM5O1rFxexbSwUVrhKB8=
`protect END_PROTECTED
