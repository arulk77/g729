`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42mPfZva5hN/i4nQEtBzfNwIX1+Bp6wOY0XBmfVKa6yb
HW+B2KUMGe/yIDaQxrMWLup99/r0NS0KCPxsMtSPKknnX3yePr2CFFkahug51qWh
TEPYywUewdtJ4JC/aN63uw9+/Z4AvUc+RtafsTPSEEAEaCk3KbBUCZfWJlBX66ng
CAv13qPqnYktJ3fDUc+MTHV1Int3zKd/ormEVz6a3tHad4/1R5kDJNEA9jNo84jc
/O0OFIHmMkIkPOE5/w1m5WPpLN08DvV6j4kq7CQzM+2yaw1FnN7uT4r1fYWvoKxR
nf9u81p7L92i8OvszVPe3w==
`protect END_PROTECTED
