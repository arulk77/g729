`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eju63lrAseGy08hZA9im4YBYKIjcu/OafZ38KxplGgHKBA0dQDXJXfAgtAhl3r8Z
XLF81xjVZM538Zo0lHue+RhUb6KeDukzeLYdJsZjcZCb7vvO0euYfC1Ns85Y5y1j
sXkelelycWS0bm2d8ro97Q624VFlvaV9bECQBGbXkfIAOn8ewhCx27dO+KArBr3E
DdEjtV1YqvCDntFB0A7qWCFIcTieUueNrMBzyhCVGWgXDW4V4pm/xGiKFnUGMj+U
fwAtkPF1wZvrd68BRP4ZQDQtOx2mDtGOjnXcIbFY6gMC7w3VmOHEELO+aUPAP9mB
4WV0nNNk4QftnOCW8PJD96hnxtgk8cboJDQZz+hgNd5S3XlOf1JJBMiVW3jWFlUx
vLN9b/kfhT++2BspADPu+n1TgLdf8cWPmVSfx0DyUQxBWE6fpNTEVhSCiSZfArFr
JxCSMwBjvIRz05Kh3uzTjkCopMHha+8TFzlhryoULZ3ocHnKHuTqQGZ7pXQFhBv2
FXMdU5HnjHzce/6bScd9gkDXVaHZ+mjE8QIU1rrUSDC0zpwp2UdkEP8onN3KLEYs
+hzpyQBpvtM/NX9QBgDJtg==
`protect END_PROTECTED
