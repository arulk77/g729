`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGMkjj6YOghTbModq+lbP15BcJrhfnPld7giV/AXX58k
xCl/Ke4+TPS4in57gb2ywB8UMsV+jHhWwzx7x4I0fRg2E7vGPHy/W2v3lLD92Zxq
0oKbot3T3C/DbtwNpzTBIpkj4aFsVOSu8Rii21QEHi3YoE3oPr9W8jwJ4xybJRyN
uWkqA4mmjfvbIkt8Ru44RWJ6TNa3SKWlONCNYxAV6vLTPpjJi4mj6+QqZauac/wB
oU4leRYu6PYn4igiBL0QvNC6yfNFvmADNY/BL3McslbCAfzdJgvsjIcDTbgYH0Kh
Y0K8bR1xS4tZsagsSGSBp+JpPhKLQwF9fcL1Gvixlo5PZ8S+MI57bfZepZSDz7pV
qKPaokTQrw3n+xDikDd1fOB2aKSONxt66xtnspZBq2waGWSTLKM5NwnNgYBthm4n
STKb75cILh1+W3DgUxxVPHfnpMrNZgo82cX7KCSFxhWedSs7JmzqYNHSYHi0iU09
pouv/b3bny6++wrboMaJEtEOJ0H/jZoEuWXmue56cVJySc8gAFAqN8JaQcppl1c5
JuVt1mcT2w8KRPbLoHfn8/SrLg0KC0z0/oE28gO86qHnyevfJncjji6UPZsoNLaM
jusOz0wcVE8cvR5pJB4NquNcuu4pGFIcVFGRrtctJlD1FFYQVMW6gWUNutoICMgG
lyP8iY+sOWIuOTzI0OZYKwGinekfWMdst4JW09OE0nfEM7gWI9m5px5lKgZ1rO8i
pxICedryLh9ImEFslZGcTbj98IRNWfYS8B5K6vnrx4+OzmJm2rSPz0dV9M25gCQg
/r0cInTiaqQ2liaH8+lkFGMPJVT17v5+5E9L9vIHmFij9VjhzOfNnZARynHsXTHl
gScLa4dQgM6GX9N9xXJk+805vpaiVkHsf6Mw/UA9phkoYwoliOiVf8fWu2/ecb+t
Xur0rMb/LMyYxynVNgBqrHgHr8+ntQBKAEUrkQmECfVTs4grufQMe3rV+HoCiSZJ
xRbFoJxe9VYVU6kyKXhaU/NClf46V6omL3HpfuzDq1x46uh4CnBn6cRwOIJyODCf
SntszzYVOKf1ZvUvzXNKbMc8WpNFlRQXiuiv5e8+Ijt0NdX/1CoAL2VYBIOXmYqZ
ps+lOAYUthIWIjJQgUMZRZdXdn5KD3cRdgVHfJx0b8chkAoVeokxsIaf4WElsFRP
vNjt3hj8se8GnFZx6wtjvSXJD6OziRF8nHPCgwQYVdRY7N09vCBZ6R++qKjnJ2fS
LtHoBp9CEpPgoFssJvFlzN49R+TKuNysoJcthDOtNg2GFjyaBhLU8FaAzX3lBcXk
A3+/d5/2E3sNDPXfTP1hpq0oX2q+79QThLZ2PgsCnSs+LwZTBKy+POwAWga1kv+L
avGW4xjvwYGItpQOktnx4gKN3yOsFnMvyMiQLG76NtS4vkPE5Vko/zlNqBK839lL
8J/bfJKo/PlE7H+k01/XD/PNQDl1L/v29S7o59WOnVhYXqyVk8qmN6+wcy4Rseti
9+/yESRil4rGFddzrEMloQ==
`protect END_PROTECTED
