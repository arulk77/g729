`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePJlQsX43/UmwXO36+OTnDnn7MiHgLN8q4cYqooM7HZn
PkJ4LBhzYYvV+vJUtFAvsILKJG1b11SRYRIZA4s3osMiWMR6p4UFDwjblErVCvnF
oGn8dxlXukk8ym+JLtZw/G+GAQ+phkDOl9vMrUcTOB9xehfOwUGva5+TQOUBMG2I
QLyLHwNKaxmj9bw3niXMB+mXDAxUmQrowU31Ck1JxfeeuIMHvoJ51dREdTm9deMg
`protect END_PROTECTED
