`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mTKd2p5sd6hsxuvJff8fakDibtFAhB1UfO5BQe06ohnwGzhqvQKhNqhTpwaUga1j
UnfFOpZPIZDJVQbWo66a5CCI3MCmukKCPrrxCsPC+o0tAZ+G9odxjUnnLCuh+doe
DEsjHF1TJpsWm9sIgDCla1EmJa+z/KkTRxvV7IdzDEp1VCZnSMfyBXKX7PVnLonW
TvtB1eNjWrg0jJQEA9oTNzMCjC7Ens6iIIDZMFikPrw=
`protect END_PROTECTED
