`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEGerJx+kASsKAPRlbowbhfd/f0xa2c8uA9/QaR/d5ib
R54SlqxlICBsvHvVqNQWyI9J9LBOpF61vIbnNeRY49R1FLB3gPyuPAhMMX5Ewr1H
/CTuF9eFPyWJq2jcWs/oG4TFC6ZbVoH1qjjm+645aXYaCQoqzSOpeQbUoyuOvDCQ
xwlx8U5fDuVNyO7/8rG1070g1MnRoGEh5KDQ4Mgukx6nKCGgzJqS5ajnhoNelpsn
y2XbMMe/NPPBI3Wk2PJKC88HHJCM8ijXzGfhQ55MGyQul4EydTJ3oZb2w0ql0ql7
FW5uoIME1hGCSdk6VwJui9iD9jYWv+vYB09coMm8WgXCNpT0YFlfORHmhoTFszmc
CN1KlMWZZpcA1YVHFZ93xg==
`protect END_PROTECTED
