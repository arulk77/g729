`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9EbHISG+boUo6thuMD9rHR7UzDX0xAMvKQketFKIjTqOtsh5mJlsM9eHPUVShT53
O4XQLfcHY7+vv59FBVokawnBCf50vN58nA/lm/InrfMY6haOm+fxZKlXYiu0ADB6
7tYzynPllGAolRSfkYAdVa96o8COipECS140cssMOuY05ppj3TjyEUYOy21Mqo5+
JOPjDReIeSBNYaOoQTixBG+bclDQ10Vk5nDmW0MnBkEjjfhJtryiMKeGVFbZh5cm
zlPUcJPy89/gvp/XDVNLHi9C4wx3N+FkqWeq93hTZT6yshJdXNB+4SwURpO5+7rz
pk4ZdIN8ZlmpaAEFpXY9o9OYzVO0REi3QzhARH7lCeho2a82I22kmiXBFKT2hGjq
lS4MwV+ULqS3rHB4fgUjmGuqbStGrDE0oFNEqY04qu3MUtmaVyc+pNspsviY+6QT
JeiHCpICF6H3rKCLKW6VZlPQnsOeaGEgbuscRQuism9R3Zdv5W8/dfujKfGhQPhF
bd1WurC3z749TwF40a4DHf8UwNt8nH1Hr7hqj7q9EPibwJmOT6O1Zo01pjoHjMiW
0lnsrC0oQYBMxYcNPcUH2aBYdK36gfMMnIz5qxMXtihU/DS60D26yG9J6Jspc6E1
My1xcwfLuKMjMi03Ub78w6fIEKSpz3/xp2FB2UpcKq9Leoh1SA/qoZn9Z/X3JsLv
pZPy8p3+vbbcWLt9CnYTpfnDzZTj3Vrf96EC2bfKlb58tf5nx+8kjWuZ2s43SOVk
CsqpGfK0LPuPYjiEPOxTnYlvyLSD0zUVsRilQLm6ajqs+NlJehsn7VtkIFzv3nvj
G3OD2x8F9gGK0UFYjOiCQd6qViuhP0RZ7Ic/WDje12DmBSlC8MYYggSGQqHzXoSO
B99ov7Cn5ad5noV1vmzDBdeOCQoKvQlaEstBkAXIZ+BlU3PwoKLX1vgH/a8ahTli
A1ufU4Of4C7ysH6Xrm+TuUYnJY59vRTjX7cq47sf57vitgTo12/ZvHOXwopLDjv/
BbbFVecMuoZOJ6LW9e5a5ApEw/bPVEFauEpcdjws1BbdwIVWOl6G5xfyh5lh+K9W
3ORHyg3F5o4GSngGeUipk9CzADqyMr1a1p5nZpZILbAOic+4pPd0vjIHCpwGK3m8
tsJUp5g6jpjgVDm6PjMdjv8WfTxBo4P4URSyeYg2T1Bhp3UAQva4a8hXS3Dsbs2t
b+YvnYvXs9BMV70h54sXH9ThhQpUZxIBiu7pHlBpV8RffUD4qT+wBVpU5j3RKpm1
7F7Tmpe2IdydleM8naed4I47mo7IIRnjdkKjHS8rY9o26i7FWTEnyOdHeGSqOk+Y
wrxU3v/lkgOcOb/wVtNU96WEBAYPEhNAAYYVVq4xvLzG2Yr0CkRcNq1P4DRYQREW
wqjnyGC8kXUjALRjN4CH26S+5mlk3G1w/qlfxnEMrfo0nJ11xezA5QISfEOYD9cI
WfGXKL1m3Jzn78XysTOLHwRaPcaejWAk6E8ssGfMdCN19s8xgkzeGcCRo1cGKNGe
5dr/BzYlxeyoziAiOv7bCx2m0JUagj8W/abl29IttgNacCW3hL+2kZJUDH3LuN0m
baT9Z6rILru6xLQrbNB1WIl9LbMaLkEDlkhc8cwZ7kh5+iTGiBHsFvrzWUEBouw0
cXjKmA9uXKQ4V6jk+wLN9YB3ZvL0rANqRTirLW70gRx59fqkcautSgJM0hdPfFoN
g/XBw8O2MhlH/JjEc1pVk6vLVBNpO+Z9flM1dVxoQ5hCFpTuw/g5tqnXjt8MrT3z
xFkS21HN/fj/KSsXElgBZkeIpzwWnL55c01qI1isIh/OcF2aa+bQRkw5RpNgBPxD
H47LUh4B8d5RB6ivmu8/nlLECUTasPlPkkhlsAToTT/9WdYPz6aNGJdEYMoO6IXZ
lslqQfwp0GoSSOe2A8wHrylZHKaSg8Wzl3dnRI7aoaN9XUznxe2KHA36y2M9OPaJ
mSITYxLbvR1EB2XZrfCMLA4W3OzAD/EXP/LZMx+TovOv1y4Gk6W4neB4gHdRVFox
NMXwXzfh7HWFak/3VJPHPVT2Jr7Kzr2BYqHGic6TYkiw2tj+OlfPnrEYx2gVe1T3
GOBtQNZi0ZzoDLRtJgOCPdrvcoStKmbGKD8XfmIraMP9WGjGBB2TVHRk12HOqYDb
YY8jvN7KfiXd11LJ6td7F6eiLik0yeS7l3/yjM3QMLHvIKgvR6K21vRw+QYKFI8r
Ej4WTiYiswvyCRPFQ4CM0El8AuCMGvRFZDb7KGSaqutJZ48llImW8E1Iw/oXMjlb
ilQjh26YlwGPyL2K6wj7whYoaMJ4DxdgV6gBRio/Wpz25IwLAXA4OUrxMLMRSnQd
ADu1MEHY1e8Mlj2ZAdqgHqx1MHKVnuXJnDuDEYa394mapu2qIYrIKnXtGBFj+CdN
tBmRnxt5PzOoaZ7V8sdxe2BfmE5pHU7GafHBHwCQu3tkWLtjxu88W9dS0loJsq9a
K1mHIGAR4IRySNdea0gAguDSu41EVmNORkoeRwYH4hxMLBo53sIrZUy3CAItu8Co
flXSW7zGEyR436NoyAIpFpFDfHSNqiVLeMgoAcHpzHCFgeGw9+qQYJFNBoL+HklI
kNgQth0FYbExe7irpXi90hmmyQOKfwORbnQtGSRzHCfei6j08rAWiRmjhGp9c7ZR
IlpqAoaeS7SvVzOiBCQLzJUr2sTH9YqZU4AVQeZ3mnrXmsUUAiTGVLw5T+LqEpcL
CI+CabXyN3GjNeugAO9T0/9zcK9JZNf7Z3DWVo0/Bjv/VgyzbI+yK78Lp040xafa
swHz/xj8ImEm+6aqrHigAMu99VIJQZKniu+zFVx2lfrCH00oDMd2Y6FAInBTZ9hV
CxafdgbIaGsMgoZ6pN3TVGPsemjL1dxaTLMYZrZQCyO7d0wqOxPVfy3k0pwBMMuk
gwG4GDJILSvv+J2Cy7IfwnZJWPKiF235DqHv0NmQ5H6G6NiBSJZZDMigJPmcpyvw
j9eHdVNWvE4n54qxMbduvKDRKgE2XbwulKXSUYCoPUnyZ2zMmHYYX0y9zHJDJMsP
6yafKt/0pILxCio0KQ0L2amDAmq4csElzh9wPLupN4TIl2hzmN/dsx8hKvmm4hBb
+RIFDRJ/VMjlVp8iUHWX9z6BXAMoSfhGK1q6Ps+e+4IVWWrGPKqhx/GheyToVyxR
43p6UzuGVh+6qt0dKAFmDqWvwR3H82IzZoyWJQorH6hiG/eBPsB1z/VyuTE4+j1T
eReKoDz6sD+K3UCJy24EWKtWx0NKmwNQrergs0TJDdcbHfvlbV3mVOzH/xgmUCPJ
in0Df3OP5Qa1bbbuZXMcq8GMSyGRS/HARQLrmrdOsz0nyR+VM0HqyA0K3zBxz2qF
htFT8WYFX/alGxZDzi0uZcdIbg2X5Ve/U80inxwwblsPBLRdkMF4QcjJdEjDemDx
IFpbdwmBRGtSfAYhHf3dPwwYh3I4jLX/P+YywsjCM8ZhngByO97abLp1lgY0tKT+
CQa8qAUyqe5efm+cID6iH3OJ8eJImxdj3b5QyXCR/hYd8PjgR/ymXtIruAPq8Pf4
4NG+G0abpnP96iPe8WZ8+jnXoHCW3jPEKrBhEL3Sqb/uer98fSgVZyv8omy6WWgg
Z/D5vwDeIyj+HcjpeDMggG28HaywU3fxIT7iZ/uYzgnnVB0awtWkSywfDQL4iZet
xE9FREWHaTaN29ziD437nI6//2e2Bcze7JOF5uoUV+4tik+lHMDpqRFxzJWnp0pk
tNbF9mM2Wrw1a0GUNawVTrphjpx391EsFoOo7l2TcQCNkjjBtQ66hcsbLh3gpRZy
S8gI4r0qRX3Re6eaT6S5H7eqJB5PVdhXb6PKB9EHGS8ILMTj2uYbP81I6L7sGr80
SQckvGqgSyPKkvyNbmlafZfKv2zL+gYJrFFn3EQ+Lt/WHP0271QfUN2U482brIQ+
wX4YJo0I2WBPeYvW8HAdsOlhUZDjGVFMWXNcbduxJW7VITS5d1VBjCRUHj263vKw
RdmJBLxE3a6MP1XymgoDTtrCJaC4I4RwJ+NrBmMjclBL9CahVripGjqiX87kbbta
PlI9GdnVWYua/zr4zjtjfpOR6E8kX1C+sK/lAj/9cekLPnVJbPpxxbdfamKtAh+Q
2JuLqWrEFkiIGODolsBKv3CpPgtNYlIk/2MzrM9l8Jinq/DWdtmUjRW7oVVlMUvA
ES0PunhDSF5JTc4GhByzVei1koXh6UuTkAtcf+sBva8CnbZOcnMnYbYXc5+9UIHF
WSSC1VSd6nwjeWpwaBB+Cjlzn4dlDMejDK6VgDRcyhUNjYoIwh8MKtpNiiCGfZJo
hdcULmWsH2cd//SRfaQ0+VNTTKqappkQKQqK+JU7SaYtgLRmI1lWNv0HkmKWO1F0
i9qUFJbDCwgVrWCujlPLwkmBSbiy8LVtCShfRBqteVLT6YtuFgByz6d4f5hIYLyU
zqZvfedGChDRKG3qRJp0A+4crHHZxmVnj4iMwIwaDAfvT1sgmUt3NPPIfUfKo3V4
yCBCM3SbtrEXIyrDZ5/UeTGar3u8aTt14Qy6gts1VatNPp7pRhUHWmkXV5uPNi/M
RkDHPFswW3jDXKUdxMBZXIqVGVprfE4owlBu5NASG4WEgmeoLD6APxt/SaveBMXu
DkgW+qpo1u17yo1+KkPPNcS1BN0kzQSlfdqB60dM3snV6+4iDtITCELPXFNnVTZi
itS9BoOhWr4gW/tgp46VKu4uV10LgT006VsqBen/hwl0ki0W9hZNbXM1LMo9THb4
u46cV3TY74zpTzMkK5trS5Gf1Rz2WDmCj74dEGfcDnc10GYvBYB47LYAkrqOk4fI
ZbuJIcbPq8crTxBuWVFoHE2M0kmYeYN0pGZmSl5t7og8QpZyMXhOz/sNJV8Sj+tl
3ho7MckUyovNQH/K+l4Pc+tstls/2+3moNRncrZa6MvqqDNpKBc2ArkC/r93N3wi
acnpLTyqrFXpEtKzhRu/lA/1ydUnEWnMRYcBaDy5Mz+65za0/sOiXkFxtp/xhQWw
2q3qHQDPIcr+F0QzLsWflPWdc7JgfnzZkWnnuboTEbFzT7XacIvZ1sWnSl5zJXvT
/rop6tkgxWA3oIn8bbGcinj6aFoCqt/AnMS0zRrQzZ6cBUq7ydQHQ3v/R8vBazfg
bc3gtYIiR55EX9rnH+1boOCSBN75dKK3CiS0H9PaWaw9iEF7TEVNL3UhOFsQQydR
0YzNQP59mmq6yn/kJYOr6KSSli930np3dg+8LSYJrEL/1z8EzjntXHbZysBY8zpz
vOSCC+R/8z5krvv3Fd8rlQTkbW8YokrRYK5HcJRo2g6S+t+XORn2TTm91F7i/sE5
kWJv6liq9RZ/U08oX9/uwB/Qmfyfqqzj8E/Ysx8gqSvAdTf+0PIssItpWT8yihq5
keNIS6u+s7IBvPQniTbKfpSwTdxFrX9+FDj2/Akwk79Dy6WjtmTG8LnAiE3ennLz
B/sL6BXxqlY2bbxa2nikLP9uzbBZ18oFuAEXmQGMv3H9wsYeSzNQsWFIK0qV141c
mINX3+0vrRBIuWl2cR2IsdGDiheyUmEEPXs07PUBbso+TjaUrGtyt2CL9GIkd0gJ
FD0SO4ZRIuaYV9PjRVSyE9GQWlU4blpHvWLAxqAy0rgJFsxSl4b/cpbX20SjVwQE
gm1pWyG2jz2BziFujgWJdVvS98dgukoteMTg7uFKMuaD+hkHr2ixiA65FtVDV+Vz
LndiESQn2/awxiMK7zev2NlOp2fbF3reYWsLUuLePJ/JQ4McPh2pIX2WK1BUbrHe
nQ/slztHau+R26/HQtorm8w1oN2nSCTwBb/NkTYxJnGP9bpqGSTC/wrTC4dueRjX
RjSos4+gB/6E62dB64Tqb0de+XTtNxkbnLhC7pLOCtoFtZosdnubBVUaXM83RoBT
7qYaBS0BpttZD8rumUljr6CxecCIW9e3kH3Ia68KYiOoAfhX81FsvjlHDqTszO6R
nHV+UAzdMrbcaXnhHC5+Zjz6BHS9F3WYABJknWTS7l9HYXsG6KV/camVsITGwTiQ
ecxNq5y+nJ5hqjHz61XMa+wB/nqqRr0RhG/HwmBY0X0nm7tEA9IBZy9tD1k/DJKD
t3LlmD0uPLsNHW0KDgcwAm3TG2NiQz6hFZYMVSzkrqohtRhHtW0JJU6x9Lc0ntWQ
kQOxi94O5TvybZ6yp6AtW3ZV04wqZ+9EzPI5gE3y9dNtFfFVlD23SxlVqRGAFz8i
yFdUfN0cvi1coH5+geG8cnWLNE/3HGVyyedb5G3Zd5UUfg1PYZW0UXFnOtCHarRV
HuGuBJi/aRK8KbfvhCwvDJD+uYulvaaPogJjfzZf2le20jySnCa5POog+IELg1G2
NVB5ODynHmtB0GNhlfWIMhJXjJccURI+rAoY9z42qst2tm0avF/Sf0CrG5Kly3Ln
oSTRV9PV6FYB9ICgY0jbIpQ4rO1DVpzIbzmv/OZdE4o/KR4Ewo4DjtIYT2HJSJY1
0dI6J6TMdO1kZDTDevAuOxBXy/Gxf4NmWOUf9UT5CbJvNjcIrs3z1W7ioXAG+oCy
fI7FHiDMNfeIeNo+A4I5yl6WNKYX2gltjIXDKBnDauCkGAujqA+kvfqYXbpxtYKx
BI4a5oN3JEBXIKcR0TkpdiKyo/9qdlRQGp1wuek0+h3QP3K1SNiUVXA9vK3DVNQu
5ACqgcZ4IqyIAUku8iJYnINxcak6w7/DXHC9iUXLDAUG/BcHIcvnO0+XAr7OMCyF
tFC9vLySGTfLYDA6ApqrkSEzUnKAXIxRU3UcFfg9BcWGfR3suXJUZNh2IzWhb9LK
mGtLC0fweJXGnzHvf61sd7a2jdr4gqEWuomentEU8c7x+TqgMVIH64yUpYuzeafI
AfqVAkYTks2c38KvKVesn5xG+CpqCwZpJKpRRBoZmWihJgC7jHrs/hyny0dEd0ht
m4FU2JA4pcQ5mdmASAyYc7crUcfic1vrJs0qSPp4SIrfyhWRRIXPon3uSfPh+fKB
pp5v+ef9MoFwWcqd7Xxpk/qYzgzadssw7CutofGBe4W3fygQkUvwjBodO9J0lny1
EA13x9gJwBH12gC4NI1gUyVKPaA5s/ZyZigpNurqDT7zVaJ9y08/TAQj92X1d5kL
5jdBFxfgOHNeW5ugh6PrAPs1U909qrNSXE1lHs8CvCxzPo/T8/fHqyLQAclBHAwF
5+qqJCYZ7PuNjbhXmLmFCBOvw0z/tnmVo6LJGWCm9EoDHLXO+sC17cKCmuSBajx3
sQXleOtvFOG4jVfpM59n6fJN7K/+uqpFw3aTV3d2OauEtVdPgmzprbMrh95WZrRd
te8+lTJNwPGrraORHPWHZImolIsgt8JRVYKNA0YJ68mktRNSaZI4w91wNbJnPerf
koRxWB5+v+I5WS3rfm/BVuTcAFllXyY8VxM2TFMgrmstuKYEc+Du7UXnbrhkFVWs
UGMca1seYXv809RxdAh0dCVSQD275cv7qUqx4Wi6hTn/05Hug4NB39gRg+XN34zF
PYEb7vOR7T1MYrnDanZoOLf3yLxNw/E7ijM8/CgTiZP8Stnfy6/aJTrzPj9tJncp
tz3wbfeV8ew4Nb2E4YhDkzoplhWZefsvrm+PYYeZRWxjqk4rSFC4+12VI8LCY/W/
RcDVkpre3yY+C5P669PXTQNtEta4TbFN/L4TJaWEnfuZ+DJCB/M4HqskVXkuV5kR
lYGoFjPFrMMg+dDLJpzMzYXVak1BFnsqKCGUam4Psd7tLtr4molLj0SimCaM5x31
/DDBF+UI1Bj58xMsrDT8DcKUCU2RPLKB7q0HEzqBjk7GFpq/r4cdSZ7PQk8rJLcL
zZsUbPmR/KVhuRVyV9v8rp9wA763KwHXXJKYCGP8XTPf37iez1a28no8KNNjsehD
EKu7JquLpa5+9VB2jnJcRK9IYYBOBj85yBmWeyn0UN6bqR/dyf1BAeoCqPjvXdID
6yKIqoxbKS7kCPrsn2un5JizJ8Xkm8BOEvgDddSIv2lj5DcR6OM1p1k0m9DlG4ZU
8bKmq4MalGkTVhNAf+j2AK7r06KlmbQhlkmT+HSV4h3nXJju59StTbb+2SveuV2t
6ONWUX0yiPnAwe3r35nywODSJ1Q3DDSYFVLm16YtaMlRga0H24Q04WbJC5qoWqFv
qETVYpTPP3gIjfBwhs0DlyRbL9f6Om5/TmHVo8qz0pPFiOGk1KX6+V0qcsdKUdPA
jVeFQRoBRqyTI85h+EklBnH5VIeK8noUdqzSQDbgFil5wo5dSgy2GZRTusrdl1NX
IBWG2VToQ3uFTkYq+gMEuREN5zyWvhWfqLCfGWonDikyYN/9Y9S0jcKRj53nbYuV
PGFi9VMQIMi4K4kccNCzakDpLNa26TfRm0jFf9QpWVDFpKv24va+lnefbFnuig2s
9grNKQNakrWpxtgJnXdTh9tr7XgqEg7/4MJequU6/4+yw2T5ZuWatEu3mBvLSydj
aPdFhSlbu1k2jHO3NIWzAVA6xJFlgYpjW1qNopjeLrPr8FzWslYsd/WDWqKckUyX
ZqOwGuLICrzvj5knWE8v5y6/57VA74ZrUq7CaE/b817vwjbWUpFrqFBv/nrEinJC
yJoDuHjzQ7bvOH+C4xwyFHZpKXq8lXkhNyAz5Nu1z7D2rgZEFC07VTjTAWsnKXAF
/BKFtUDSRzyPZaC781gAw+6jqONeCO58ZaOSTF77WDIDGldh8EjqGEYJ8loT6/IS
lvqjRWbNcm3YXFU6tNyKDd3hZlU+zb0dmsUXr/hFBZaXCcgqlboFLHuVC2H053En
vXno3t9vD6cLROSmqqcT/OAh7oXe89HCDhGSfr8msEp7e8JdWQVEDpDk1GZb3ZSD
AvcZI2qeeW5ESVmal1RovfTj4+SQQojmFecVs+hpmMDaiZG3f1ITP27r0u15KxZN
ocqXFhvBB86Ccl9fOI+h1pnyeRdqKeE4BwYq9kHFcT9DhD/g4BErjQtEBGaCw+50
UqonF5OFrxIFaanRr6eRG3pY/kgLEXLucJ/gvma2Z51E2VcPh/cw7upDWCx1Y7GH
xJs3ABQdUBd3BOQQX9c9/+u+cUdo98kbRFXNwV1dRqsgVEhuEt7niSZsdp0xEprG
kl3dfj8JE217ibczqW7i+rfOi/J/YfJyKrIvsPB06C6m+eHJM9ay2pUkcKPDybPl
55WENWrTzrtp+lLmNUhc8nq05Fbo/mbiFrTJfFo0yFVCcmDgBKrc+ljCMBHws8+x
mrOb41T1PKMdalDSmOsnaI3Z1SfSLOT12Eqj9YKA0ueWtaTJndjcUpVrrFgdAOTr
e7Vui2U7J72/UcnH6MOk5RsEsZ/tqVpOrHeudNaPoDPOx7k5ebyQxDWMMli/me8j
f35yeicU2nqoYqmQpHDFlOuY4r2Ktux8VTAmStBpKIVHdjw+LUDIyA8fDcX7Z9fP
1pVmiEAdE9/bulVjDuBAjV2qWyzOHBeu2H3temPQEOxLnWpDUo/tnj4gt1gSWGng
ty05KPZZpwgqmuh55MKBVLTSF2CNtWn/is81ZR+C3XY6d2r6p8OI02LfH6qmjRwx
OAElKjxi2qPesRzjhAXn9JYNM2+PQqrQKkGLuGzF7wHaZurEqlELPTIqos15qFJx
x+k2rUNNzZm1SR8zb26TkxKnL/s/vOtylBFF9CuKhAHYvKP3d3Sjkpi3QLE04WvF
/MVLiU5IGa7Y6DlzHmk4WIJKG1x4skpQKf8L7nchJaHPE7hKMiW6J+bk3HL7OdmM
lgQd6SNO2Zkyz7ICvPAgmQhIFEhUIR5frj4/gT0r9rLaBHGxPENgNSB3ISOIxlpT
BLOoNKBkQOqOJbVydVbHnr7VR8k2Ir5xgt9jEpSZByJSX+dpUAxJrt5BwCNUfyGw
Gi1dA0S4zjkxky53JcOAmQ+prvyw1/IhITkbTvOiOAdqrMQoRq/uoS7DQwUAu4dl
FF0WSG4pfnPhfKmz3AObcPPJDVHotvkBdAK609TGw8yj/h13SuhB/1nIMOOK96u6
NX2c3rhuW1vi6KV17FN7jt/THSso2Qa6yFkTbv4lwGwy13kXPQQSjOUytQg1MGK4
9esLPUAmUwuW05PbhAdMigz95zLpi5CR7sOPfBlUT0uHStC0pRJhAnGFfu01gfwd
6zi+nmT32YvDkHVKyhd9HzrO9bOHy7yDLpb/YYeqDu9Ugt3mFy/UumPsnoVgJ3UN
Ea20nOanzDDeVPNbU6y7xK284ALglV+1GT0FC9cIfdUQ6tAiHBRWH62i07iDkRiE
GqBAp0lQPNJ2kR7EIGYiSZEgOydXl3JcYMbIRRTAWkPRHnIIXso/pTFAkFqIqw/0
aFTpv2ngAzyNrWj2SioaQT1BLlqrxWHJt6tL6l81lZZevFmQ6OwgyQqJL6r8f7hK
Nfu2wVJNQ+XWIxZxj07nJypqucM2OGk44R7+gTbVg97n4PVV/nfTOzeAIatrz96h
A2WN2QYVCCsUtmsQ2gWKNoG1GU3lqsfKwvOhQ97XInTYTSdqY3tE4kyNKE3zEW9K
mGXY6AB30xMKo8eUH5DyE0IdTAweSmQn8kmfmqI/PMLSFDFM4syHEg332IZfMamT
o3B855Zk0gqbdUumrFV+6jA4x2oatQeHTKZbWG8EtaCw8lXHc+RwaEhqNxjILj73
rUt2Hu2ZM+ZwnPcEw0yoBhaY6nqB+Nr8Xtcj5t1s1/hqJ3zte93N17VMFUzoIpRp
/vRzr518Ex35wQovw1LNleJz4jpxwdoJsuEKJ1rL/kO7hGkrX016Ra2mCa8CWJtI
/BAEti35A2yKnlRWR3DAz2MHTkovioSIVbK6Cpg3lUFqeVrCv3SL6mbONRenckBX
q+QhPofqU5uPLDdyAR+7EL2qK9o+SDRJBgwsXxroIm0SYr09KwOkoXgOrIw+8xA3
Gr5FJURhvYMIO0ocCcLmfmhU5nIuxA2+ytZqmkNBjg1EVKCyBrTr5NgtuhoFIPk/
xlKeZpZOBVmXu2j+/+nMGxnhvTBFkjrkh6fWNwfePAQOZlOqH6tcWq8DTbZwDYet
tl+TDXuPWodHsZnVXw4QM9ADIlOOvLKlCdZ1ukjdGgNyI6ZEMvdqfHqKZnE9pXX1
CO9N65wAenDl0U7PbkG5+xTfu4iWAHT49kQOmvhsqIPZ4SCvNjWOKfPf8MrPhVSL
TGFTP2aKGfo1+Op3apUpbmfqoX+FcWyFpKgFGrUIZJi/+VNa0XPPcYruBLoDqZMI
bbEqDmCP/3KoKi5xdeGloIogUZzWDxMXHpUWC/d9f6Az5HuIwsNt4N20gXN5HaGI
BDvVrTLvmCKj9MIzU7++dXNxxAlY6X+VEJiOpeCaChGTNOcs0LVvepdQGCJpiBdc
D1bh6WD1ipG1TAozdPrOSg8MBE02Sfg0hU1AAh5wvS0dNHaF7hFaVR4wXO8tcmow
HeMatwUeH9TXidmqMEMlMrmoEQPMSSmgeZw3hnzzMcl4E64acgYWE3zd1SrYo5UV
g+J6T/SFcsFN3wc1B79V7qfcKjrZBdHv2sMuzD5X5dBrRsES+gKUSert+qWMo26A
ZUUOPJitzrM4/E3dIvHLFP0ZpltVVDuHYypp6Ib8C3iJplsDuEsiSVsG6NO+AI4K
yKYNsSsxUPwq+Mn54GaAD+pib5yi+IM3/Vb0qzRLP/53wbbRnnxIXrHrf6K3RPnV
Fzo3y5c2Qn+mll6XP2DKC/49WQfo6qSzKt2eoR4Ou9G4rrvXzd4o8kBgoV06mjb5
uNfNgYPzJr78mQHZV9TouT9xbqfybe5lg1rgQciHJzjRsP7KcXSbbS+6VRRrBSjC
bji69G7FROOZ4+cHUwq97Z6ZpkBGPphr+xAXtD0TROM2pJs3XjM2qR5hhTMvo5fK
raGgLh4o8oVAzH2N7OQYRTPjz5TBSxcY2UUkRGiee6knFI0b6TAw2xwRNxO8beC5
tZKs2lC5WdmvrACTeFavFcC7yUjuz5hzAlYiELnu8y9HQPoOcTegKqnZ3ZhDT10X
6y/T+bGyTopS+qD8m7zQrY7zAbyAZjZ5r3XfOjolUfpFzgH/XQmhnb/fpMWR1I5B
chVg0DiCGNziCLsb5M79kb22IUOoamAPMcZlgcqdujBMebRI864ZRuz63YFbbIfx
mVWMdq+1W1rRek8fwa6NJn6Gs+GdwIaRCRfexd0y/wW3ZZMTZEiQwJmhBjaxqyXJ
lHAFmmE1KvNgcb/V6A7syRljPXe1p81k2tURXOSFBn2aUmp+s9KwlJYXKZr0taJW
U9f+U15WGr4F4W19ivG8klSPdH949Po+DLRr2Oj6B6V+Mrw/Ks+KZWu6BhhF3x6p
+D9k323y4BJCGBe8R9+IDYyOpQRuyJ77qLxCH9YWFx5KIFoZ67cgPPY7jbh4v9k7
tsm3gL+mnT+2QDm5RIJa64yW2tyITPJp9uYFUjxODA+yjM4cz0oeHGFL0ABSsHyg
X+12ZkytD7ERE1338kAaqzOuNByn+iqqGEXSqYGObhGO9ep9zMhuxaq3G+1gjyDs
3O91zwrpmL7mhntt7KFN/sQ/5mwgXUsRJw+XvZzWPlMYMm30yGgSYtLfp6t7ypgn
ktp4CxNHyMvshVFXkRoQ3iMLY7RhZiWXT/hLeXO0w+5NcKDV3N6+mEb77HafZLWu
tDqQPW2ceALMEhSVjTQbRYAe8MhRNw0sOnKto5fTLHJCDWzMXClZo2K62Ieiovgg
cfLwHTjq/oYzXvdFjw4dUNDzg1L6DcbcJZ3M7zh2d/9p7UN6QDn80IWCENTe5KHr
wmw3x3b1zWe2tzSMgafAZdV2K1oilFBZ604Tibff+740XIyjyjVurFO6s5yuBnz+
2DTrdqW38+PueAMugexTifgY5f95SqAZv40mhJb+/7PBc1Iw2U2YTJDSZUDXem7w
Ud2CThUJyxc/5/wJdn2DdLDbXUsv0hWYyk+hMGjTsq8hugB9eJf+n1oip0dcfkMc
0Grc9wheM0j3h9juZeqFVb306mQzc41pwE0yeKAgAZDItqg9/lN5nqchOWtEgxc2
/T+a3LxOXZ7LwKSmPNd5HQZdbuFm55dHH3V1+dmDBRLnlooc/8rCz+HWe/PECi6v
M0MixN8ClLLB4rQYnbXU54xzb6+9z1EZg8Kcz8KNiOyxtAbZJAvSbEzarSKWYPfr
Hefm4Hi8Sxm538vu633AB0OzYwtRum9b8FbQ2LsQiEWlc8ruDH8yv0gFgFS/7GlU
t8by+ioZ5bIM/UNb2POaHKNgZTAwI9vz6sKiaYSzaiBNKa8DF00CbyOHjzmBClGA
rBxNV8j/MibkQ9OyqFc1yqOCaKpvQpLmk+7VccGS2/PnkSHTIjJ5DBNs6cBpZriR
TIvIPTysj0bQZUCS+Xf4UtL64hh/3WeMUvGGCkL76Ie8BI5zV6aEUSp16WRvryWj
gZ9G1BJli8ouMFBbam7sFVkzRXrREUn5i9/DNh94lrqJYs+CoWFDo49Syfg6rOAy
qldw8dYVHfyX6Oyl9at3aqZOpaHn2RPadVWroTrJE/5FD4LgFc0A1D1MxIUSEXuP
hIw/oB670pHaf34LlsaLuNmFNpuuXqJOhCMq/a7ciXx0nl+cpYPvSh5pZekDYjhE
Inp2O4GHkAVa9yh8KyvZNk4jRzo5Xx9zGOHOQK5iNikUHohhPwGq/yt7+AwJ6V2r
ur8+K2FRZ55+PCkRnIAoaOcEyTZ+og1OLF6nhOPxjvrRCuNMn5dcscP1icZJSWbW
hDoTNxtGEYSonQs7/qx3CsjE/5te8keVpaPxvvx3ANuaxzD4ZV6o5bQQYWON4qgV
OiAbj1m6umIrUQY7mZOutp19b+TcLQPjPZH9fi8Tu7kwcifjqC0TFIbItz3rnsZB
0gXHOAcyd7Qi0FUC/4DHzJPnBN2FpbfAonSWQu42mP7+ZCyzVITue1B8Dwqgr3EX
bfsSGe54C5DN6xNVj07JvW6ByC67xE2DHiusz7cP0pezw2y4ZLxFCLmlTjrdHRDC
mdrd8hOM5k+stujNvtEA4FJcbW8pU65GcMxVPczjkhaWbWVXUQS/AGoRpd8B/kWc
CI3zwH/rwPvhyajIHSijDpE1OfiZ5dZnMbCl9VGMpY9+3iGLikbMD1nThubFnU6l
VfoKp2uRGlkyc+YCWbRY/4UbEJcJL/1sMjMSJgig/cF6bLU/nTglZcOHJHEtT+qi
LUrhcltDo/YO58LA3CZzm89IPvEifPGZqzexFQmULyGnDIO0E/MoeCH9M430SKzU
zIafFmJdfuWYeF5ZRNyfYVnijoL4KIkwmzrwYjvy3jH7qO4Mw6gzr4OyNdze0I6a
aJwwLi1rZVQWhNylu1GU8OfWR63USo4jOWBGpyH90Nqjy8ATUSPLqm6AAYESBgMv
e9Cw1LbUS5O9g7B2DltsBuAmzqJa9/hLIBuOqtSBkUSwQ+BOcLl3YPSSy1sJlAJc
SYyB1LHrL40tKO7PQFjKdyq0Hs27v9ouPQjVVbsbrI5/HgtuH1tKBjRj2CNwb/fg
BuqR3mu2CFqFrBcNKyT8a9j/WHa4PYEAoks5n+R4D6h+NdOF72TznIjg0/XOI/DO
+mqeq9j99AhVGZmsSFoXD9loHOQu9NtNUVm0A162TXBQoMWtz6gGpnqdUmF1L6P+
nGVsjYbepC0nIEndhA+j9SJF9iXd9w2hxISc/8GxdYeB8ZvrUmpf2qyC0WwMf++s
JX/Jkp7yK0x6hgQFZ+wVfOVooL/WFdEtSB6RdY0rhm4lwWPGBbCRHsuM3aF11IhD
JbB3Wuxq2Ryjmj2AcF1SVwF+JLCHafbtj2153Wej1lqm0DjML1/1S6oyqRSnAMAn
EpBLbvE5tACKqieCu5sHV2GP3g4FvgqP1hqnKJzqY+XG3ovYdF3kKkFh9LFNmq9z
3NGgqFMBltUavPCIsFopZfBqDXuZxSzXroZftYMZ1lXe4XtM/7lCsGgy+xmNYJq6
0p4wflumdEqsxv1sAfNsTRw+SqUCN3LjZm0hmZw7K6/HrVez8iYaRJu9gEZ/8e63
uZEDKX0ZO9lYySwEuT9uFYDMHRxEv/nOyOw8rjetqa7aSETLL+hylVlSc+t+JxWS
0JGQz38Ocakw4EKxIum9tahM/CTadSWDQLl71wzBj5/q01+JoEIYr7yJXn8PmUdF
kZ4rNkkV8i7U+HyNxGCBThfJNWfmdVK6gykBd7nWMF5OTrjL2/41+w6a9YhXu/nn
ZRkT9h/7IYDJfAmF1o6ZGUurU/jvHK9lqN1X5pdYvc5YLpdwtuwBkg7b347bbxM9
7YO5Kh/0JnZSfhv8pqrxGBBbaGKICyEhemiJj/sxPhZp42/HCSjSwaorpPMoTBFT
8TXQg3nDXReegZNFsTHxRyb+YL01VPnoUZBpv+W1UYvKgvIlVjf/zL8hWGuNeWCq
6u1+9wc3NSjyQPrB5H2I5L5gGUHlWaPtI4UIzZX4sTC56NYxr5wum0It8CMQqUzv
ZOU7D0IUTZQq+Fw/FL303aqa/GLEMWuB3CcllN71OdsyEwcHqnI9j8YRGFcMMS6q
8D+h8+Pa2tFq9mfcslxU5jPiGgc4Ab/0pDhOQ6g8zO1HtvRIM3/c9qkRGRTxLD7l
oc9scvfVARWgJs+YC0BPqK3V4jlQRRagPCECYv3eaZgdW5M7UtACqsNF/7FOTgke
/l7dZopWw3QeXk9UnnSO2jsnmFiodTjEVucFh+vvjc+4sXFXZLaMYccyBFwAmJom
2K/GA0NPukzWlyTO5jRDh/X7cECXJaw2Jw1963ODErxNKM3Jxfx0RtTvSpZPPxIy
9QJs5EDBmOkWAc7+fnZUBxEBuQVEF4MKF1QKF2nnCgKiHMPbU4fQ7KSh+JbkqdDu
kf10fxQN/LmgCeL0nj89Nmm8snzN5mC6PVU9wSXum/Nh8359//y+Yw9jI8Snlc3y
vdJ8EGplFMU5RlMGIW4BVONHuU4TpTsl+qorv1Nwgb3MqQfMlKBK8sWJjpKy8t2V
v/6crWMEdYVKGvyYBumvPl+x7zY8VruEBlEa1fNi4kB5sOgDri/ap4CcNpNaiJkj
ujMWwbai01P6ymmgIbFxQmyUzNlDwOjkflXqtbP4HQWlE8d7TDxcZ7HwCEBTTAyW
cabNdEavQkx2J+qjv8ImXhPyjuUfG3khhX0T5bzo7qhqMs0vncYelx1bPlvx5Z0Z
kxGkttDStpPNTaRCqiOY6cNm2fC3aJ+trt9syLBaalXRnbRtrw+62BJxFlk3PlZA
uo5CGnXC6d1gioRi2YS8gTtrnAO1SchBJmnNpnCdADT430jQVQhV3Aw51Zfe8wXT
z8XaUY0FwXPjR0ddqb+B9DgxFQHzb2cj19xeBaxDgx9VWYeF922yAY657IDiVmP5
TeQGFXql98xAmDBi16mQtnzgdtff/je3vigpKH95hYKYobgPghgpa7oqPRxP6La6
Jf8nbI9RB7z1KytiEAKmZT7TAyJkr/TzczyCBzg6Ci4beug238VrYOLrN1uBGtip
718uvSqLKTFmLjO584rwP+w3aL8lPW9VvlvrzsXxeJeVgmgHqRZRz1P9M2CyMRHb
pe09yURCNMrwptMLNAbeF8AbQ3wOdvVRNYGrFwPvTLPYD927zs/CISe3oaxa7S/X
HwAb8QSjkHefpUEuDPJ2a6RKEZ8qP/q7cIL1CQBpo2cdH3H2oVw7PdJ9Ajr189kI
lJ+MHXkY7beMAiypNRlV/EpHed5k0xxajBwZLIGTm/L7SSwalz0VE+QQaNzkAMbv
tXbwshLfpgxSxcDIWwpRef9dZcIZbaqTW6DWK20/biWDld6jB29xI0wpnzskyFUB
zqDnUDMJtfsTss+7oFP99JOkRnhDOh5cRmmSBAKzNc/i7U8OSqEjYODv0B1QEOoF
++8X9DI0vv6/Lf8E5Z588x5M+5t2PjcGq3gbtB+uruahz01pfDJKQZmb0+UmKJs/
gWMjaO8lAfHgRJDr46uEjSVPZrpNWnnpHh00z53avsQXNImNqaQAbJgW1S9RMH7C
4SaLalWCZDPRePEKhHMgZRduewGNiYp1G+nyJFS4rL2xchQPbam2UzfGsRKb23wk
j2XES/nA3knPESssNMIQe4Aw9AeMgfrCewzCcWqZjuI=
`protect END_PROTECTED
