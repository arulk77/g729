`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHqa14kwI/HBAxMZ2o8T3kVcwUIyUyoHxXpOejaV6BBq
4fbFFajEFFuakbiDDtEPurIl2xVaOI+H3aSRr6Pyl05fybni3XUtiyFK8UAt25Fl
Q0ROWN0vfUw6ABfgXKxvXpZ7tgiSpzDL2gsNmqOEXZJMO51ZxM5lDuOJnALCTPyd
xUFzhXQr+aEk4UN6XQmo7zLOR+kXfDxxrT2F2MLCwLCrc+Soi4l7I6QwSj+UymOB
MejA2+TopkDp9UbfCF8iSP+I+6flzc8y2hWN/GTsYz16evFP6Ub4Ygj6aGR+rNm4
SHuI/L0ONTMSJnYgj0A9PRWomS6Q9Mb4ZftZHJaUEFoMj7/SH+woANbijSjbeUaM
uhNLb+mWvJTmhSZEF7zguoOZbwnb42xOnzFQmxPlUP1prlqnZzLX8HrNNqaEb++0
zbNYbBG1VSJEGGyfK8X6LPVMnlmw7to5/8bMFfobq8Fkon4onJ+ltPDY9BHaImkX
U4ANHAKFg7YtyI+BQozh9b4hi87tvU3vc4avtr9BvIfPiUXOGPMFyhI+L0w4odwu
`protect END_PROTECTED
