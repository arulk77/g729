`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76gQczUFxxV81HCRH7tjXkZFNcEbmFDkjV8lTWKkEcfV4mQeIq9ZEe0eHUf+S4rM
dGoq9sZB2iMrx2VtOdqaO05bjyvHdrlHrFKki9p1Oayh+tThmG9IH5odGfMeNcmO
zrAB7FYcqpZYt8f29gmpXUmgIT3PDU8O6uZgyoAiHlBkhykZvvKFDO8hP29WZXbK
3Lpi06AZ+ESE9p4IQpsZP3kcbL/f8R/TfXvPeRo9BCb+Y1fBFWKZA5Fl+6BuybUE
`protect END_PROTECTED
