`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFAMWTesaxmqitAxs/jUS1k+5wKvGtyXv48ddQGuMFuW
SS08E+9BXTT7yvGtl155M+OL6rY53se1EcjQQ6Aq2uglhtKtCtHs1IMukHH8eR+a
clwss8lKBnTruDWptcbsxmFEpM8cbbzWaVwd2hx3rx9xTJJV1iowRi/FlFp6zvVk
X1hY1gHw4iCoKehs06MJWdF/2R0iaZb/1khq25dAluokz6Q2u7oRXilTTWB7UGB0
IJhkVOVQcUqM0H5uQc7U7w==
`protect END_PROTECTED
