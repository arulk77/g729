`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SRQRsRGBT/BOcqGJi/lh2wDHZ0IplDLC0r0XcUPoKMRC
iS/AIgF3NSchhp1pYB348/eqf/0H5rK8yuWnXfzRcbiyddWi+QC49h76tD8+3PrJ
urfx4zGn3E2RL44PaFXeRvuxiulbvaqGnpJAYlaQ9ABNumS12BWBBenqbE57XC50
3wVnV/Dc/nyjPKcxC64a339oGb9DVlxcKYP204765ikvUsqCS4yEHvmYdnaGhFiv
7jkSSU6TOb+SkhXWgvJmGLrOdCcb5xnsyw/95e1hYKsIZDS/OJ6DaSPBaBcy+swn
/Rwx6dYcXe6KUsxCXnfC+g==
`protect END_PROTECTED
