`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rzh/tPE6Iv5fglWsZF7uo2DycYpCsPyrPX4nuanDs96/rd8PfRT1wWfX0qHTp+fT
naB6vAi6+nmqwH1xhkn++y1TTnQz4kF7+g5ja2ljv/tuD3wr959RE73GJB0lDl3m
pcd6NX1WvM8QIZWX2Wn8h51VLqeGWIQt2TzvXqt7IR6L7d3eaDDczhvGLS6gMk9I
sZ86zgleVVhoYE547wE9bxWr7h12r+ruTorIu+qHiF4jfLeR7+bLC3vk8KwBqbpI
dxOnPSP/oyVUv3doSHslfU9rma//tBKL7J3F3V9TDcWumLzXpXjoNVKafMoFBwdw
dSaAZOHVaCT2tPMpq/jyskXo3Jn0Uv2oZThVLmp0Hq3U5CxlRXH0ZNIj+36fDg1o
FNUzAVvXvIHlkB96+b9/qmXJyfLa4Be6tERVKEEGVMcfTGHSP8te2NzSRGxbVpDR
Ibo/iVVh9zmiEQdkUhwaar4MzQ8ZFvuxy/faaliDIaFAKAVlHmyouCmKE50lnxj9
L+zuHZ61b7Lo5qbJ1p9SrUDnVTthSk0wTB7uf4t276G6GXUEqc7+XErg0Zxh4lbn
e7KaVLr5JJCZT/0Urf9CBil3N6AuInL2V/VWzd2ZpsJNJ1YGBjXpAR3l6wZroFCv
S6gf3Zn4sUG3G6xvgeSo19NYkyei4QasDpHCTcrKJ/xhDlvHpgcRAvviE7D8INnQ
hz6HQU4CZPVrjO3V/xMMCXefUAuvLpF0LBzURWQ3ntlyMkFJtWNLUBhnn6KrGVVd
S5A8kon8hejtA/pOp+YOzvqBRMpMzFjzQYSDmgR7lK+dbA8V+K6pnuxb8dQSfl7L
uN/QthtJonNMcWHJ2SrMlNan8hXqdSIO4mb74e8OztNQkv+41Qw8V6QTUezfMyf7
uSWloAL+6fxjhQ3CH683Wlxv29HSYknFaH6QsE9fuhRzl72wvR/H1gfGnV65R8af
CDbwcG6T2p76rR+COJ37/SbJTja8u+/Uk7hw7mY9cOH7270gKKxgli9C3/myp/+f
OZdTDDWzpE1B2+Tkxf+36S2reTpc4EDI/0DSVTvXkNPdhLDf2M6CblaHWkxrlWM7
kRp6oZl7NDSEfAQHBzPqoKGNPGl+mkavZE6Z8uY+udStAObT9+nQxZ0EkkOQ6CA4
2UG1gcWCxEa0iis3GhC6OxJqssWo9ikEa9pq8kyH9Q9+kW6u7n4oZ9dWzBmPTPSK
OrRWgZZX8wZKHsuZ+zUL38KE07ZmfpR5gssd6CnvpO3tVKZYrnlk+nxcclNTLggL
DnesGNkfZ28RsWeA/oFxVq05v/vaA8dP2P6HTyXzJ8iOv00cQuMguWashTZGS9Em
D8O1yZWckkEApjb4D2V6aBIhlD0MG3bsX8qUryh90rnkt9RwFLe9oGNj3kdGGCPZ
31AIyu0ByHUGjrjXR0WnSfOvxpAcy9nz38wMbBpPK/EWRSfJHHIsgujURIUcVgBk
5VibmuhJhRj6M25HK8LX6gNOjwVv3k6kNHzcIYPO3uG0mXUCGx2uYe7a0SFdgPve
nrg0g9/Z97qlz4aJ0VUKNk9KaMpQXOrLzKyuQ9/v4MOsmlvueEmVEEjpFBRpfALy
o8Lm54ETP2F7Dk21T5TUTMQEaYbI/TPTHPNuZ5EWwdGvSCZa5QOHe+9QZNsPuZtn
2u8kW4KItTyPnZghNfqA2gPlAvtuFgmw5DFJIdlJiFWPFlhv70rHZ4CJ+RuFHZTU
4/Jt1fmEnJzvxqxwvNk+MNNWYeMs40YDQCUfj/y/C7hMKW6i18nljoygybRNiwAG
0piBpX/480zcOSf/2gvn3xr4wTAzcOq1TZ66tol/YIHLlc8vVQwsbQxxDbFUZHcu
mrsjQo9lGIyrddKiHUuzzIzS9ZV/HheBkOnzfZhN9ktp7nZykZWQ2ej61zUhbif8
qdFdeiHhUAlsInSyz47VowVeTGwt0TATMEjAC696fZNDKnS1sqktkPdLkMdY7UyD
NItj8VnnVAwB0NLpPNL2NP7NllKtO7TxGQ9bNFQoC1UjHusju/aI3M1XCCnS9UHB
9kU3/pZ4IsTyB3ofHz5Pnr5VmcOvzkq4JKhxbTsBADBjyVZhbfo2jzMK+YjjKpbR
IE+5BG8DQG3FmIBhdAOlCFHqGuFvRHr7TY30ZarkB/02zI52d5ECf+radvj+yy+G
j28n2ylgKhz3Jrbe6mfqPkNHEyBcup/HMiuFcn4feowbQC4fHpDiZZdrAien2eQw
kbYEZfWljIjGd+poGUq0qjbh7/MRtm1OmrYe27leuIhtx5L5t1OSPcDBrsP1MSpA
meoFYoamNukYMc4cTeLdXSfy7EmjnNCatWqichvPcGlcvrpiDeiFmDcmgk5H3T28
le6iENc8tgEa//igZyJOJw==
`protect END_PROTECTED
