`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE1S8cnH6DMnKK0Vc2AWHDqV3ZyCOOlIXdmmbNBACivV
rWOxFwYBNVzcpHWKag9OijY/vkdVzcHrthLBiUAOpV8w2W9qMuTZesFGlvWBbM6S
l+uap6KamVP7sq3B5rdzwawBGL7NT+xzKUnqmBpsweAS1h7CTzJ4en9ZVxB5sA5v
1ryekorZzUcQeUIJTeWjW3JrK921NnOA1OLuKHkoRkZ7qBGLncLWO94Ck7o1NlD3
`protect END_PROTECTED
