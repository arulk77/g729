`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xktFbQ9qdL32ne6ljkrO3XJ7tmWjmexlAKhuyhjkkt5
YdXfxpKA3OBXsltM61DTamuELujgOsMPT0g5oT+TSITBw/iQwFF72S1K0O7iZ8nM
ZirhupWZqxdokNORcH0chCslhA62IRHka9ARSKac38C/WHeKRqQE+u+FRTDruDbz
WGF2diPfLEd/iwIrqkiyoVFhrXqWVjAU8f4HkzlIT2vRhRARhlVAR6jjoNjXPFqT
1wJyvI1Vk/uE/H+Lnrrmycsd5N02O6ZrfT+emxlXBoc=
`protect END_PROTECTED
