`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI5wDChJYX8LGUbLJXKcqQ+lhvYUjql1YPAT5r9WX15p
J6RwdYMMMvCuTchP3yNjymNJUE2iy6BGrMkYRVcz7zC0yhqWUoME1SWW8aACAi8Z
koGuz4lpY0DyL3liSm49nLCuZmzRRWQ+XMiDUNhi8IfOxK877LmnzeTZVdFR+bUK
swYLcoLjC/DqQRBTOcCTpBoR3UnYEShWy1TnsbPbBa4=
`protect END_PROTECTED
