`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43C4Bk22ZkFm6CjFyWeJQQS4/2pthYNQI7JYSiT8M6zB
w5050l17kIoOEH4knIBnVavgeNIxWpokZwmhWyw58MFXmwnb17EZQqIs1IBGBtG+
PyQRbR8jtMoArnSfB3hGMLRFlXH/louYmBvuFcLhA2MHdwWfzqiQfFdg3Cwj280F
GJARTau4ZG2szUAMFZOMH8aZncPdDWVMMZmzQYk6lKpZ6lKz4NeUX9uX2+kNW6x+
7G8KzlcxR+1hcCUXHU+lQEEYWFXtW9upvP8aW2tOg7Pph7AW2nR2HR/eNCOKracE
LeUBGFsIi4UiGF0i/tu+iQ==
`protect END_PROTECTED
