`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UuKKg99AC7RPKIo0YgDm4gXFBvquqFAI4sXCLBXwVCE5zJ8bqgwXazLMloBvCvH8
ET+DdH/KwWVEc3Ocm4XwT3iM5sQzhW63ANUTTPptfUEvPh8QRU+XuV8ti18WaJIX
MaUhfMw/gHnKC1lLuVtzDCokv80dpTbp0eV23PQt48xkPpFbAni8udW0vbePR2RE
JkljvhX43NgA0vRhT8opRZ/kV8nhl2EzdhcjlLpzHzOz9eJzvwFckQmTQ7R4Sz8d
v2kqcIp+sPVKzRMuCpP+G1FOxtZE26+wn+vIxvbhdY/qdqZGZR7FL2T18P0Yniuh
ph7TolEmckxcm5IxrNVX+jGXQuTYjn1fi4HwrchXpZajhbcu4NuNkhZ+DniaNg6w
Oz6S5nshRM5OnKkpbaO/njC9Fgmw37ttJXsVTokNGdxMn5Yk2TR7TCaVtnEp2zyH
swKNod/JEIAqbxoe2IX5iVNp2vWhX1BNkKxmA7gzAmdnqlS7YzmySjE+/36yPj3/
ZT/a0hLoZhzqmRmuR5AdcN4xJX3Ku1HxcTIopTUk3zpMaFMlSlXjl95GH+oownBL
PqRYsCmukoL9QHwjc9NlAg==
`protect END_PROTECTED
