`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOkknNCgHB8XFVeXgM6b40sXCs+dHQwaXOtARtGitgK5
yUW1Zt8wugnjb5cXPkROgsNkvapnteYzcTqh4MlG1K22ecYgp+M2zIdrbLuPtlvm
9gaYgejrMXt161vcg12kS4nlcZg+O2l+remptaIE1fMCqITLfegrBtl/CFtC6gKz
4BXAfYue3YSWOV+4hSjCCg==
`protect END_PROTECTED
