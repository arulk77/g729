`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN+GGlwlCk/fLYNXbaBsXBbu1Tfev01qVIGZqK+lQuTw8
6B5efGvVdVAmxoBF6Aa54Nr+CTl5wbg4nRyQmOu9M+H0+icJ1y/fVcdeim0FjGJc
1l/qenUuOZCW9rk2lodZxxYjY/C8ByTy02CRXY6iBm4LdDy5tcZ0t1YmwH3SOExz
9ZfPf6B/PBfb8GCDYSJ2PdsenQDXTjhY8Ryp/AcTlhjEZhsMNiZfVL8gv44VyyxZ
QBp5B4ItbXvspxpuI8pp5/Oq0cZE54ihuh5hgMXRn1yM4WHRx7uIXkQbzDDRiEzw
VRZvzGq1TiZPffgiHrsru6TmZbGfhYYHWrpYdHLKIwR+oThB0GvR4L3eEiswu1mT
h60f1jLTZ+dNd5D8uqg6H3fTTHkzkXgHLmpOpAl0Ikp3k5tT+5BBMU+CoUFebIWo
hvbEhewA51rSbiEziwpsKPniMF8OLumka9fpDIIYg62g/aC570C2hvTK+rCIk3H0
0KQJqNZuc/9+kYAYCJC8wMuh/QJLlIvBHRpdbPGtKMFnqj/TYG/LDAJ1F14d0+kY
dud+mr0T8K5HSUmPIzoWTmcU08i6TlEp6wTgxdu+xIVgrTjJktk6xL4pXaHek2dz
L7H60FLzvGm7l9D/2Trc+clGDFCkbjaLIOdALyXYMZ5M/prWa5Z8pGd91GaizQCY
g/x0cVd+qT1+2EUlzY90NHnrUTBVtlU7aly+y4GIRSgL/J8Fj77uijjAUtjI+zed
/DsSvswcBtqSzmib/dzO68Enexh4yi3hhmO1+6AE4v9gMGskYb5qgtmTUcnHVk79
EHyCj2ck7VmaSNTeRwij+kWe7faNmT3sA1VOS8nGcf9ZwpZEWU5DYuaeWjhZrzbR
cs6wHOek2ayfpXnyG3GiGBkVL6SQMtps6h05NrncXWt23f6ULDaPvoihPM711xG/
ncovAZka9PH6qRfvqKN0WRV3ifkrH1B6660RhoN05brQ0Zs1KLFQ2Jrf6/cLcGpU
UujvmXkPO3EFfKTmTi7gJ3nrLe6ggVJPw1BbjwPbEKQtttt9ISucAY6udc9vjT/r
aJxxKi9az6K1oYBn4tB8Fjar7rwOqqrtsAWY70lPBs/ZrCN/5OkIHXlT+Pk4dPIA
2fVgME0u5gh9dTQ9r9OhVDIR4aOC7RN9H20q7fH4My3ja3E2PlKzijV+nbzXKf/z
GAIucCwj9GB1a3E9SGYIpA==
`protect END_PROTECTED
