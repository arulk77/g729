`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQNY8/9SEfIzB71zce7sODZiX3AzsnhtEZ46MqvHFGO4
nyQ0QiN/xJ6WrrJ/9Wv/wlHAvX28W1I/UUff5Wc+NlLLkHPLgnvzLTBPP+W1d+oE
jMzZ9d7TUyMDIE5X+cx0S8XfNmh2noDA0Ix3qEDD89KlSsfZBFrVXNYAPOpD0D9F
czuknQR41DmgekuhnUgdMa69itlST/GgYn8UfIL3B0ayDfFrhlaE5EvS8GKABAez
ETpRiUTjq9h/4KSETxcpiXXMdaF8euR+W5My89QFee0yQHeoHqP8v87MPqcDRpzh
6+I9do0hl5UkKYkfm6o33oLZd37Q/DeX2pviwV3SbONGfqEnjTQeHmW4lS/AZ2qy
lIurMWGJVuME6wy4y++0oBZ/gdrr6/dLGjuCZs4hbhVZ5GaF0dr9pcJzL0z6kN1o
Ndqj+QmzIUtI+dePlkiRQPgQ2tO9XthCpOy5HqWDvgkS+q0dhtcYHk1gibHnwMni
ukesfcx49KrnC34eXZSDW6Zni+j/Lnvlv4ZkBRi9KRKL2LonVxrjuWFGpEGakvom
2iDD2rROmW8/mTYH2swZ0zp1XZSSCdKGHnGFVBS4MYY=
`protect END_PROTECTED
