`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zVTLQXLurHfWhLhicNhCGZ2tvW0erlcn3XWamAeE8Qj
hzQM7b1C9bojSByk+l3jtNEN5gKZ4Y7Tzi34yceN3hfqNrxUzHyPSdQJ+Cf2hToI
S8jfptQzlGooBoOJTZttrwHwyjk8j4Qp9xfEj1p9T808pQYkYGL7vgBZd8uxRBHD
FLcDGAgtqWa5XaXNEyETHJusaAGmQvAHQvBzL3eAMrass8q86it0vqzQsE86VbEo
/DPf81sL1ZzrGJvsACLdKfUiBUbS2csDmhWILiE7+sU=
`protect END_PROTECTED
