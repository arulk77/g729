`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QM8fL9rzo2R2BFNZVLrb+prNAk/+L5q+/k4S6bizTZ6pARIkGwJZgMdgJxWotRcv
7eVCmqpt5IIkOB1Bc57N7R9IvtVzpcJsLJJxv+opcyZjO/tYLvTxqvDOV9AD5wAi
`protect END_PROTECTED
