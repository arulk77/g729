`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+8ZCZmaLnLHbmXAIygKgV3g/1CzSDKn5/zaNVrIp1WH
73/BxUZTCIyjSTO3HisPXrldHVbWATXS6+4VdXjVMpAXNfwqboYH5umVkOJMJYXz
nsnzour+ISd1Nuuoj1Md+NqD7bg+0nuzPTCU74HRRwiMibZTLOXhG71GxY1vPpV7
kgmibGM9ugkIeV0IVozppPOkf/puz1iH8yp+hBFlykjHdwdHNzJtKt1+jgl/heaL
ccWc97bfFN8d3KQCQZJaNozXB1LgZU1TDwoLVK5zlXxCSnQhl2sxZboqfnbbNUfS
tG9fHpjiccZc97LUhyhsBfoYzz8xVhIPsouOXFP9r/6S9ER4i3juLms0wydjfeUw
Ut84SYSYBLkCtxkNHsOD+4lzDOdCZUgCQJZZv1uLruKaMmMH5RVEXKi/yQhlAO1L
KJdQLVlyTRe/4RuQvJBNTYJPHeJh5GXXI3ei5mMgACWi+Re2+11ukamAV+mzGN8S
NJrnadcrquovsltIxAMLEw==
`protect END_PROTECTED
