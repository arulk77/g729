`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMOogapaqlkdRmXrEVyEZfhsL+pKIqBr5wmmCiERTY9p
i4KPyDWQ8I+PpK6Fj5eT/oADY66fx+4GO9PE8jtF+wlGqu3WtyLxSWXIhhcbVB7i
GwzCkUyfbdSNVtvYwufeCdYm31YWe/9/4p7HbGRdOp6tLrcFCbRrz7fY7xpss4Km
temmPjE0iQFEs0W03x78mds/tn69KxjDoeHvolzFeEGkaWL1WKDXMOw/hSixYc/C
gJD6uMEgLoePvx8SPQ3f6CPEPVgbGhjunIX1iPZhg2qybRbYldcR3elXyUf0pzHJ
3YERGC+cnTucF+kD9SVkrBuuwJdUJC32Hwe9mwN2LLIDxvCmtCtZwoKeRlUZJpvu
RzrKB85hqKnG7vDVLKnsyPXPim89ESHL4s494FHwohhSzfmI3SqKeM6zrfHUoObC
SqlGdNu93qebh/Gd75zKgxWQykbteh+D+DbIFgjy5HB2QcUKtBlKVM/QeYM6AcRL
TkKTltnWCAtNnKiQTXJoow==
`protect END_PROTECTED
