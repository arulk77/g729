`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA9GMbP/e3P2i18Lgn2a4tSI5j2oBWdQvpC7RaptSxDs
dp0nWUClpoqqxRrQ9jhK4lyXEqAKGhzvc5YPedkWxDIBa07Q5OWHGPWhV0/fQz2g
XZzSaYDTeFq2Cj/veIJ8ybpU4dmMnb4MbTTAo6sKYdtP1/1Z0dxy2/isGqJ+od3L
zn02cAh9wasVDOU5DBXKDQ==
`protect END_PROTECTED
