`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN5BMctS3Lu/6zkMlf/l0bUXQhBShfmDoAJALGYw73ht
WjVHu7RGw9LA2nH/dkhWy2Ewn3cjqNzIcIxjG2al1p8qy8CjPNsBbyukg/Vh2l0t
NOGLaFpQqvhOFR5q+fJQQSn4KGXcaSk9RPr+q6wSv3g7uI4iNk84G4PYudmZP4cy
mON1OSPFF0f5b3Vw4uJ517v8uB6aKtgpx3bLOmHQLVJBY3VN+S0WGj7MGmZyOGPw
JxECdBzpguA7Iq5B8B86d1mcH+ZGwUWZA5aWsKuE3nOkLsubfTbDlsVsloCg7mwJ
DPs/OCTNl6VH3aqquDxLso5iyBmspl8xCCYWWKHQiYFmsTKfknR660AZe/Mz1sG9
XqB48VIXe4OmRjfNX/06gCMx4ZUnSCdNJYtEbfgIa0qWxISSCn7BhNgCL4SbZTgg
5Q00ZmIeApd3BqGmf3s0lSg8BijswGWZ2oztmwsqF9mROYzjR4kK6jZDbL/gdNfV
SNgo4+z3JtpfDnwDmmgEHpQZpnVTaN1AvU5PrCEIsPvlWOXCkUJXnPo+Q6gA+egC
1/7TQSJJH6BBqgvte+p2dg==
`protect END_PROTECTED
