`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDASOlpa1FncIPFdrK4V0JWg3E5MQROm0enT23afnuCAVz
HmFAp/bak2drdZOfQ4Jxn2fOBs+kqF1Gg4r6fKTE5Ct1ZBIxn2xZhztK2SOm3G8j
SOPy6qWgTVpEr4STAHrVuxEO/8E3Dq8NlGdtmGU7yEtsf3phki82ykZ00aj/N/kI
oAljzELkkbgXfO50z9BotZjnQGr18iE/kuy7hSLB4vXrWJYCrSD/j3VocMmXzkUX
ZralADpfwrWhuH74TdyZvGVCTTqizJ7OFfs2l+ubCowes17RHSHZcjJ1SitcLNLh
avydxm5oHgkslrR7lkbGc7W/u2pV2+o73mrtC/63BrNiGdU28IXaEDECPe+LSY6l
11IiDj21SxH1SC3uBbBB8UyRSEUgT/cv9OQ8oSlm8b/3bl6fwA98JxyGMHYRAl9Z
njO4i/GiLD8FfubWUTDV92kcTJgH70iDE8mdH6LFK2lN8agsRX4MTTU5jil/pEm4
/I/gYchysst5oRmwUh/wM7BCJOSVYLyDcQLtktiPfne2nLf12kju0E/OxtYJy2Q7
ak8iV6IAg96RAuRPiA/P4E9hiSK1RVoEVbkNeZ3z4l6QYPVQjzFLXxGVtHnlnNNt
uCT6oTPfQ2IBwV+4HbHwNzij8Ur90ZHHikuBqRrdKcIWO9Iuzmm2R0cJGbyCjlhu
Po37cIEzIg7115VNnYieH3UC5teudsIv/1prW1RAShca97M5Su9mqIP0ZzFFmVx+
6avvj6k7o87Li4eNoWQBQlRrwb0EgJD+UI3HL4o1oXra28/faAw6EXXAs+rNh48e
SeGXlsDUXDqAStme013bo5MnkfS7UDp7aut9VLKmHpA73knEO1o2YwuWITdTcgsK
ryT9xPdvq8obplaZXGZLShBt9CmBLLAJtpvAfoKIlg6TlO9qjZSQ49KSKek+PPza
jM7z+rQqP6jEKh3+HGcgpXdXXrXVjAMAaL5bnc6FTtoMBqHRETk/hb6I3qE1qN/2
/WZPoZoYX/2SgER9rExG1eiPYllFwjuqTmwKAdD1N7Wa2GsrF2baF8NKUmByRkt5
93JKF30Jr53dARES2Tg7nrRaM7VBNyPweLDNXI5i7B6KGF9sXo7OS6J+LZ7TSz7A
IPv3GrCpsRVhN9bZErBEpZHo+Qa17TdxUbpyyYwRPEOV6LhhcjQmvMixPYcGeVod
UK4czo7FYkjIMSbeN2zAA9YtMSIREDdQOpQNwYekNxUyngIRmx6fXuN+5KR0PLKx
lnUdsSEmAjU25yOMtEHT2mNux3vrKTcgtEic7NWoJiizJfzqvtK6QrPzMAjFB5nR
18SRJpsW81/X64YLSx1peA==
`protect END_PROTECTED
