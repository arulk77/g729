`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO8rf5vJwS6PVj4+4FpnfoIObHDUvcOYplvY7o3IDusm
JJlT/TLvnhXLpF/hkiLpVxQUMevX1CmZNz+JpGSw9ixg1eihMnR9cGzLZD46xk4a
xEomPWxtq2IAUdZjmus2kJ2SlSrZtE9G10R9m7jy8z89KlodLMLsGj/QXb5ECfkJ
TlqLCUwwj8V7qFQZpkUME0IHet9cy4xoqviisfGzLQP+UoFRSkFSRrvkJ10aktnK
dxSFa8AsN9vhWef2oRwssY6VjsXjZZiVOQ4LbkD6QLYnr5I0sGa5kGRXrSqlhtUz
nP0J6FreCKtJFs9KHDmoWyAoY1ihjSS03RZ+qaIQkkSLIiegRW5Mfw+YQQ6+wmWA
IZpa2R2cTGkCkzUBdHip3GxxqzMptm0kiByb9ikLk4mMrMM+qFDyznOgHMYuQmfT
RHt3kQEOwPMET618FSL/TvpWlSfg28aXDnBqditRQ8WocHlYK65NaHGx95WuOV9m
7KGzFtJ2uMvurSfMQDEyg+Euza+40DcvTO1gFLeWcLzbsByLNdQ+OJX3Fom0q3ol
LMqdLFEM/RWhJGHjan63dw==
`protect END_PROTECTED
