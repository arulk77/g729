`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEW4IysMc0oOgftUCXsybYrw15L2cwUBCapmz1vIohkO
Asyl4Hg9u+gC2OOg9d37UOIeDfpuH8rSbpQTe2tEuqhSOgo1NX0QcPzCyIeC7lr2
SLL6jO7g+BHzIHExhIcPmjtajfErX+DLLhw84V7QlLtVsuRpNn7wJ9xvcCAuZFm0
TRKJtyXqehErUwjZtHwZYILfx5u7cQQe0mkbA/zdXnEp9kOBOINzqGJYjmkyAjjL
f/cabtI5oQhvXHBTBtgtnc2fijsqS9ReBOl/QIReYv4mHUOmD/knZz1o8B/cme4z
8AVEYsQwmIJ986RrLtTZF+Uh4aA4a69pbXrflHakvd9JxJwjEZ8ItXfavr5ZDZNF
tqNS3cbm1nh+W24/QuT0iqodQi9Cz0+LMB5DgoPB/V9LQD19OvkklJPeibLkaLKj
ylSmGX2lavvRDgVH5UUfpv9FUpQd9GsxceJe/8I+MJ1cEg17BcYfgEkxgS/m4IKb
U0f9pIiOZC5DHfmofjPA1vQPnHzs/ge+DqI06q0dYgMLXSTSY8A3ej3DufTYcIRj
2Of58oy81MNNVxaPSG9EKDQli4BBxELat5dZUnvS2DON4FGDrL74ddYcwSRdMve9
`protect END_PROTECTED
