`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAEchDWtTohq8J/Ocri4mzhacR7msZ5zb28UnvcKnFRx
LmlyHQqloWVQTfB5DDPqnpjlztPdH+ZttzhUUwoJ/8TRwG1gmj8DHoQOupVahN34
NGLveYQbR2H+bz5giPUPnZWfwuGppQGdnQnC/5u6pNYL7dCQn4JLzRcG0duK0Tsy
3zkKVuo8RAIxnULrP47GmQVW2DVACiTtfr63R/05Nk8tzsd/sy/YaBcgaw70syLy
`protect END_PROTECTED
