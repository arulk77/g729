`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QTRDpCJpjLAG8qTbyPtQPlZvn+GZBB9tkd7VWbwxgf3FvIR2vwML1T8/RIPA2tZT
rktDBAXnYEr8WhdxrpLICcg0ngwY8rweDumi6TA9Swh9o01yb26upi+9xEGT+tt7
1EpFW15xFrBjcJMRiK6/5d3IUgDXBAHBpmJ7KuDcwUs=
`protect END_PROTECTED
