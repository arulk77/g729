`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLcF7BmUgWxmn5dieN0NA/zstKoc6L8qNbyC9kT4ejMr
qH9W7kJvBgX3atKhRy6U9sIoHmgY2QIHlEmCo3tOf8xAKRjUcyOrm5USHMqgPLYi
PhkFYnKrgeetSye5Lo6FaJNy4dA5zL3nh0uJML4adPuy6w9G4DzkKT4gYqcxG/Y0
B0Oa0sgL3Wpq3RFY2yBlIkfEIK3ZXhhwzZfy7Kqm3wOjA4Wgs+tclh7ZBAN6+bfb
x2dG2ouSiI4I0pmmVtKas5NxFHgus5ZOmNiKHjm88Dr3royjrlCZ0Bcae6YDs006
8+p0aMuifmSpL1bRKi3cMQHO04ZGh1Sg/lqgRBW6whCFktxCwKMN2CjP/Z88ET35
FhsbwCIQOqGw3yTy4remQ+Re4I2vj5LTFGLotN4snGJu9pxpoRT74Dtr0MyGrdxn
D6pGhkfJSh1EoPzcs5C7JELGw2069c8ABGP5V6+I7vpMshF4bnOCgGG+X+NHDpvt
dHLfxk27YSzKXS3/Lh67rjfALydIrfeHUOB61XNAbd7JZPahM4xLTEachKsnZ4kL
tfPu+SzX1e04KErPexH/yKF6clk6FxOeIZvHnQ7ubTGGJyE2z7b0dHqRPLtyfFfT
46Pt6UMggF3wqORzLkGoQIS+UOirxa46wuNEx0gD+ha0IqI5cuRPQEAIIvKWa9l2
`protect END_PROTECTED
