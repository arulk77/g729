`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aeQt5FW6ZJQMBRaKkygh15piTUgeQg/q0hVZnXb9byn4
V3P+Fjqie9WrgIVVBthjmaD/5vBsGjaZx2HRYj4lQukLWL5eAK/NEwnx+Po1Y5hk
PquENxTLm+lrhofjIH/tsXsaiPjCVlNEbYog+A9brs45zyxXJHGbbD5Kg8lv6Ks7
MfPKv1vpVqpt/KyicRmAKVgM6H4Ngbk2zv007bGPhp1D5Bdth8ipDSo8h3bKKJri
UfxNqWcy0lyjrWpBJkXK3WvRjWrUMNZIC8mH6C6YxnbPZyHqMb6VmOZmtMh9Xztk
+IMGloqp9dPcza6rBCXFiyJHTFk++oAekHJm0LHKMzwe69udGR3ETwyf9KLibMxS
LANyeFIRceCBYtEs7azwN3uQfPpQ1X4Pw1+hR+MRqSRjFEceabakDs+Bsoi5qMjK
BHDsDO/ne3rQXdqiPt85xGfJQ5yMKOmNkAdpVpu7mJ9KkjR/EnSmGx/uzY0bM/0V
nBiTrH9ANPG0MDDz+YXbZIhrwnv4piTBkFPJ42hJys8LEop8YwI4laigLk2uc0dL
ibcj6Z85rzsWXvkmwR151FKzBpsFrIjRqceztNuzL5driSpJrDhTfBuwHk33vMLQ
81jnTmsvOMWx/rPV9UxNaj120/8dFNuR4pJY1525UY/scArzxVOnT7uNUeSKIrjb
wU/nadFoUQUxdB2K4m3BtiNKVMpEevSeJ/ZQVpXZcMLlWXS0qEKb48UpNPPX3ZX7
qEHTn7n8VgerBPeP74afKAhLcAm5w532ya4yQmGmur6IErL26oo66Rj/mku9+gy5
/SHz2NHjcGyFlpn83bDf5P45U6bWOHYfKOjT8D4yt20kNlcdqLvBzOMdZNAy3+90
MT8vs1zNq1EV3mmvtyz3LZZvDJQoR/Z5AJQhFPnJmVycVL2Mdvy7Mz9b/2USTD+V
1pID2LK5c/Uw+XuOj6RxKIb2OXZ0+dQLRwPwwBzZ56wjGq64yCjdsGdGXv7LwFhw
3pfaPkkbqGG2LUOMpoMgxI1kHUSqPAPqqEJZJA+/LUSZzYTstADVRA/gR90ChKkJ
QtoklmQdMBLCYdnXDI5cab51SG34urLakuqD0vhgFrrcmg2cDT900s7pLV4Hddus
kyPZyJmuxXFAcqcQNqbesw+NCJwJ1OlemiO3p6//uDS0pJoHUpkTYjWLjUFj9lBq
EYE5EiyH58ULm1sw1VA6Isroxeu1IKZ1hPJcrMCUeYBCAvZ6pj9sGMlbXreiKxj8
POSjb0i6xBJMQgJT92hMDtvqtjQAZ1UFfjzYgy4CUdA+xS1DytfNVh9BTvTVxsje
dbq9yBdvx23C+lfXx+l5h9HSQ5JRbjMyk2kk8Q1oFsZ8r4bwHEPz5/y9QvfnUJHd
lEL/tvQDyiK2aPgwcRk29yLRZziRJjg3HOUz6WMQBoejXpoEMsADahhmSdk51oPf
3SipkB+sFauQNequHxIx40/8wWAELZN3oxM0yubF5ISVfGCPI0rLA99qNPCz22Uq
we3aSCQR2Vd94ywclcMK+dBqhAiKcLO3lRZTXcSzPARLqbNGHNyjsJSbdcZoGv3M
HeMDZ1WXkFkUg81tUXtYyYdnZJraeLVgb1UugDitsZ4/F//hqGhBAV05/o0u5iDt
S0C+qvA5ppu0AosuuxVNAzHhSrJNLfpUpF58WLcZI/CqUt6oTHc7bDuoti4LdQVz
N541U9tESCQmmTgKZmrYKGjJPGa/K9uuUXn8hHt394AM2obDMisRJfw/OSIHv88f
UgT6PrMen9inh2vp5TnjT3mgvcKf66tXcia1T4V3EMYIrN568b7ZqMtx7GsaWqX8
k4koqxcalYa8DklUbJef6IJs05taP0ZZQT+VLrSuryL28OC082GO9xNqege2UCmR
aVN0PGrEk5XXUXJV712xoGGTNXqycae8ARlkg3hpV0uMzQuwmHQg8zp8ZeVqEStl
aEaQIt9ldCXcJ8boSi/PoqlhXLxnSxrajzngfcG7cxrmLBqFhzYcn5ixyCwQs/Tk
9KYZhm+NKu7JsKcu9ckf9x3deYFyNY/ce+kCKAXhLD5vgr7H3GoILlChMwUQ4qMf
bjyoWLuHGnClhSUp7Xq7C/wRUiyHPAsl6q1XOxPTwHGHTT8R4foyqDG55mVRR6ti
qrwx1fq2WxI8KHM9pBqgdoSUZjy74/k0aVSjBS4MeFgOL6PvshQ4kHmSDXQPLyw6
g75yjdd7xVLePBYpZquonoGlfoJ0eLh25sZHKKqdal5ljv28lOhEuVOOFEt+9uBV
hxcnh4GtRBSAUHsqvejP3viJUJMSKM0oFlbA/b2n7+1OdNqbuTaEFYMdfsN2r7w0
oRngaJ5JwmwsKpYpg+6LBf3qG9vI+y3koKI1R98mjrWiWOgR5qhIig/TM4PtyUjC
RLt1AHaKucI28Oec730jxCejVGNOEDQQOuT2fK4xisGCcltKrRrsDZVumFd4Oo2g
9Aj0zxm74XytIcfsyAs3UhNoiHt71nz4c5/umzMCa/7JMkhxJ7OJw5evvKhyGfPz
C6YuOMDTonWthDdjbEa15T/SB3GZ29DAkCuqui0Egx2cgRufQCCwm1+jvQFnqo6V
Ov7IaBbW0UvdIlIYb6ahvPU/gD21O6Kl56By+AsA8rV2XwYtlzfWANnlhgyKuCj/
xIKxfBBQz5XvTZDJB83mA5i8hWzuF4i3SXZVgX/At7zZICNAOyiVtbSUBTeNdEy1
bndQt449mnJll9bi1+H/nOJM/V1ey1iHEf8MnPh1Lj9j1khbl9/lJLfcutWPQiIY
7fVVxviMvKAi2QcQ3YdlTos/Tk9zxxMNd0c8aCVwbKfUBUebIdCHIIk8p5VHDl9M
c+9m7lEkGPKYQUQ+QzfrPxxJd4hl1ybJWZKS+zmU1URRaCOAcJmh+fQPK6arbXKf
vVfgTmme8z1Mt9U2wtccW2rsec+CAjSZ85RRl423TuA9C2suvjDTyCZ5a7OamOlQ
RgGSt1Tu5qjegooj5jL7mbI/m7pxZEubLH+lf94ZeEIhbDJet0kuGw8/XRpbBYZv
F6bZisT4kveyWBANrKbYxtiyMmhPywJkEu9WT0Qw9c5EykfSRevAvL3LHAC2d7RA
zVihGyc36I5Rs4y0pxA/ZMWdQLPUZvT5k+Z3B1oAS6c+3xOWqXjo91555QFP78d5
0DL73Bey9MuFSxH7QR5uyoSG8fpyNaVGsc0ggP6DCI9WToTKEzxEXNjxI3m+gu/9
hPVzHTrkfmI/n4svbSgXJYKGSFjhigA3GRtksoT+zYhqgCyRF9vdxkPIZNkj4Skk
owhlQtoIoyFz+BZDnSx1wZ3xFIdk6bvp13Ep03uQIKucZkEjwqBIIdrNJJhxv01H
kTlHuVNOpAsd/fN4hE84yRYHQX9FWH45DnM8fnRKRkhLh4ZolBYI+vhf6mzYNpCl
3UOs9Cwk9MKWf09qFNuNw17Q13OziTuiuBS83zHSFHA5jGrasKqTteSLyx3+bckm
VT/YBlcBhrGVeVHZpbcD/0VmUUZWueImcst4xEhPnETuyyDINxT4AblL62wmVX6p
voge08VdwXgX8X/h6TudMEPVFg3NqrKar7FLk13RXH/cbXwwwhTqHpt5EVjFskIf
mEx7tNg0/DzTyV9I2sx9KrE/oCtQP78bqzan2rsBM340LRi+0TObzskx/nomyFTv
rBRSQ8Jfp4QRH4/cb4qqBsqDzBYjnR/aQ9lEtQn2/SwcoEYJhN0xdg4js+Sa7B2g
PHlpFwBpgrRO4+9HlOqSE5FQfAiUsMqb0b3Mz5EVOw3ycatxL9g+ig6377KCfpfA
I4SWFzsJigz+COeuTQtNsZlepkHYSQjYHRWyPsbIrmmmOd9jOrUX5fi4rcljQm+O
1/wWGTBPSfDgfDWeqQhNXRp9PDIe137/bqbIgYY+DlzSuyOdC6FQS2LAh0mfde8d
mHODNNkLUZZSMw2eTJj/il1wCuSBmjdc4RWepWtw5gNGy1GzMUcpg1PMxLTJiipO
Fm+pXkAKlfQ5U5ysCxK1mZyChg4J5zeCrKAm+FczB922jOwZnPfId/lofkVrdveK
mptFdOhquqDeo9hEYlwNe09SZNDL+I2e2nW5PKyJncBqmt9fHY+47Iaeiv5h7amC
2KACxY3H9MPcC/MnCy7FTyHY3K6DsHDjzdJfA7HgFiPqX15dUPuHAiFc3K2Df4Dt
RrlKZDVJc1J0RdnoXYUi4xXdVWrq+CUU3Q0zx97TFpG7hWHTOjdTB5KALYREKwLm
MoXj5Kqz4+uxOEAomG0sTS8PEMxVjfE26QyKGK3emE6MbkZqHw6CL/SHFIQN5HAS
70kiwkxSDBes+VHVF62T0MkJ7kgSGCYiEOHeFpr7T5I0zh7SsXNzVt/uu2CRnELC
CJfe+DRDGYjtyvx9llIo95Gv8eDQRtZpiLtEbOUfGcqxAbCfGOTziPMlpzbruzMP
M/ifpqzNI/LM8bRHW2bIf5CR00JgI3ffP2Q5T6Mx3QCgEYPQJsJt0Ld9ogBFVWWd
u7Zim3QJ6VJ7ZGFtas6CvlX0gaHadIElLLiHRnpQduQg8yKhPy4oxxQWi8einmsh
wL8mz9UHx8fiVSrMuyxlCQ13eFhzpiS/JCFQnuPs0J467BIaienIOTirP7OdvfWC
B/ltFq7bzD1bKODizTdZ89X5mor/x4sc1v5OezadYpvRwjvWUYrww/EZo9tGvmYG
0re9x8+gGjNFb+qhJZxn10/kU3SYHCw0hpceRA0irsx0cV1PnHGd6E0DW+eaovzd
xRK2HQpfXJPOeuqqv6iT+A0s93qssuMhh/vUxScyT/ZWlbggj2/SWaoyMqMO8T1x
d8E8+I2MXPiS8y4CpP29bz7J5a69CyKzVwtoDhDG97q6cRa+MO2kq0wfkoCph/Zn
IMap4uW+oj/TEjIwRBtlsrM9D0qdfqSgtUqCsdvfEikDSADq3WOCZEKarlQoXgZt
6G4/1Gh8vrpj3ZA8fPaBtMAjVTxWbp0+p0krrdUhrjYJKxUWxE/t4MoIL8tyl1Bg
csX9p5VIcRxTaQgaLokIeTn95MxCtCfU94dxb5gQVJK1v8/FPvnW60lJA566CknH
DxKY4lignO6aiXXi6mY7xgyS7wXBbsFFNhxdUxuzDjfdfJBgeUPQuW3Z0Fkcy8Nd
PaXnd2I99WjZ0UO+VxFzgi9PXsdIhP5xvPBhRZ0MrgbLVhfaPZRH9OX9eJtJEjtU
GpHWXDhCKF8sUsAOHopmvsywbDwVNGEOkVUOGffrOgOUM1YQsvgUcnqcQec2YbR7
GImVEy9xl6gHqeyiPLhy2JZBh/rkXajD6utYc7PMrMarjoDiJ0otchKeoxlwHOrE
xPGy4K8k+612Oa4oowAZZ23bjnzp1Nruggk92qzVe4yhUTVwcYuJ09w4FV7WjVDx
AJ1683s9F7TAxAE2H07oe8H38QUsTB2zeKkZnZRdp7xFWW5Qe3cWWhXGYC9wlcYO
gKXg0LXkCN3mtOZn35ABRNrxJzubSdw4cH7a/pAYJcbMxvu8FUr4dMFEIl4koHF1
XQZ0shh+zBZumi4LOoeFl7GXLwi5njqQ3UTgKlrynjTYbjaJOtJTI2PytNvLPdWR
Sd975jmvPMshORrq0fsjgXEvcUNMU257w9hJYVR80e0n2X5q4Va7Vmcggkg8psMD
DatMILmIK0sNmQfUWFoulzmA//a3I8vq8hQqLpJYuy3vcyNtzehB81Lhj2d09Fgq
8WXnPcdUx0/dNPeNbgSeFKwtMvpoPvBNa9jtCF5/d0NPkLH6ax+hxm3QzyMShHFn
E8YpEsAOYd7xx6sMP4xHPrJ/UKSC+1DlRNObhNK59JAcNjzkrkyS8TB+ZADwm4gf
BigfYt/6fa7BeXfRyC2YoN5zKMofRU+VGMQh8kkyrFl1abwjzW/XHZn7MBatvjlA
fRzdZEUHwataxM17bUoto0sx3siA21g2RbXGlZMuILtGTWWqFzRAV9rqlJdUCJCh
6cTdBeyK8lYZsIboQtpSEWjZhsGUTBCaSZQXL6MUWQmaTKyEKVJZH9ujQlfFxX5F
UVCKk2wm0vyfwfcEMexBDTRmUwxEER0+2rhJoy5nqayeyIzkpW17nj0TqlNB56Re
RdO5qHXZM38wY7G8lZlcQFJAWbyPrEvJbNbvfzatMmIRAgdk6KBI2vol/tPuvCyp
wOh93osL0qr0p73AclpXGt9QTHosfSo9vEpEE69fsk/Q1/8EpmDpwlWnb5t0YeSL
h2XvCHHschD05GfAfZmHe0FgtTyOevx5pBFlqOutMIroQSK5VJUgntnKwCJ+Czwh
Jsy9yKjYxx6XIoZ09FSnfbrIvw8P8duOMQ0P4LmiXz5je1kSQRCTEPETwa4XD0yf
awKObyDVIUVBIWaFDXY8MThoxVjWgO1B5iyd/0Sh4661m5PZglOE6B4R54sBA/Lq
proHH9YXBAm8W991SRyvNP1VfC6EBO8ZY2k/NTzNMTMaT7RxOApKQNRP7kcYOttW
NH6xWDUeNfrx82cr5diL71AWGmgqaPNhrNlngcshh8LQQYBE2QHykNUPvyh8d2IT
QTvmNeq32S+P/6NFTzC4/rJXAt+kfr8GT6su+r+GodAxJkRB+L6UGpp5Qjr+Izoz
bQdwQIFMjgJwBxbP9nVL0b8dHu9dW8r9SYCwBJJYWh156y1i2FriIs2rPqupIIKM
ppGdZYjEYek4WfwcRxn7pNSCol3rSCV59bFJtN8cLLz8OJXt1UWkakHXxmlrkycQ
CeJzkfHem9F08IG0/LnWV7m9gBCz/hgHOYsnti8CDOEe9Nk2M9+9LRKWKk8RavvP
Kj9xMpXPGEFbQa23zbQzQWOx9mV67tBI/BKvhs6quTEJ/pHJHSVULOq4yuZXqp1h
kPKJU1TcxpDhC+cKugaFIAhOZKIWfsCpysyyETQepQM7IqrC94tlwq6btHecUh10
xmXGGJaqvXQzc2aQ/WwFfAV9ob1DpQ8sxmMJZpKZNi31fFaR/9WollE+zm0/7PvM
b3GoFwWlLepckcHBbxJXPG57Uam16S94eRMdev823lFjFB/+sYJRP4mAs+mv6eNZ
b5sJdQ64zY8XWeAcSM+9EW7gdlwduHf0/uiHkOhXdAC27nexysktcnwUMeMsQq2D
EK9KaA5+DkhVSkR+uvRDNYiv3/NDtB01VyTZYmF1a0+kjVNWp13xF9NnYUS5BIIq
dhL9OezKKIZq3GQJztg6biySdSuXC6fXeeHm7GL/2T3Dcb67+k1QyWo3vIEdKakD
yN0NvVrfwyuc+fsEKc2eiGfMwNscn3BiDv7/CT2WaTUvYbbJOY9/QwXd4ULzh4MW
TfmPQoigpIpVqVuxDCzOe4FS7fdOxq92F+0FT8IsqLRGibMtN8JfKjzfic1mz4ps
yiZAf8IP2/6ng3nae1qACR7skb+/wOsSZDiFLJLgOagCcMT4928oJMDnGAETmCb2
yhC6ADDv1ycrvnPC/o4+hwuMxS4Hzod9haDzPaLH3YIaP+y/85DZtyQoy7xAbD4c
QgHJio/cJdmvcx8KP36bN+B9eXWQgb52pVxytRATIIAe6AE4I75qKKPL8V0ObTKS
eZiSWp9XxAFRLZTdwc/+G+KADCYCRC/HYaOxFAHaOYx1ga2yEdVIxJwvj5D1hDkx
eW0jJfY2TxZLKNf8aw9stvW7gybZT1QYYRtH2QW3d55ZaiqjqNw9q961N26f9tfJ
`protect END_PROTECTED
