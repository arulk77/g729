`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C9ILTK5PrXUJFNT97hpB+DTWRuHy7mPnJuAHEUOhpsDl
FNUEL7lxUM75GmTSjVBHgB4cTzJ9Fw8Z9+WrQw3XcZFKI5Kp91ALormrfuWXk3ac
0lT/4SuHl9IUlYM/Cgje1ZrvZqYSdN/hpNPqs/ndM3UA//UbvkQtQH1aOsX/vCdm
kfhenq4axfL/UW58Wj5VcbOEWf5nFwMWwW9VB+bE23TxnPf88agx16rBBrfWb0q0
S2DfMhVSC8ZE3TWLQwLGwWhecg4qgOTYN8QyIXrelVFVF7uOyyuwAsb+hF2Y0Id5
LwD5EDkm7TAqLOFtEGStLah1HrOUiLgGbqm8XzQKoB2APYDJyc4CgE12wO+N4IGz
lNQC1q9g9GFnhs0PzuQvIw4OmKBlOvIDuPQYgWvAX+kv9SzgIy6JCrUvAhMDCNOK
nB3zKhWwiXVlxcqfH3DNgnNxW+2KbZZ4/avwrhoWDIPFiJd68gKXRRIurHO5kAiw
cSL0dBuuFhlD2X+rUHbjX8QOJXW++DX2wSvmSC3/NaDLJV3fabV7a+LEIT71EX7Q
hhTFi/Y+OrTAP8bv6OZvqBon7+oTbC1vvNwwAkfKwwDkpK+nEXWi3LiD2x+TnLn6
HqBp49snqy2XSrjmCMfLX0GqpHfyjkdCwquq955wXaAai1e4lBwU7E3kd/a3yZeQ
OzFw4LdHm3Vj9uo36HHihrRY7V5WaEQNuVD6W4zDwi1vebwy2I1xp6bzHOih6mDC
jskodSsNpWI1jkESdpCpEGMofdG0B9KvE/o8PRfZj3ThDyDV/RY7f/Ap6VqW4YPy
d8Vx0PXsuloXVqJlgI6NZVREmpRQXJtpJpo3I0Jng1F3W4jwKwO9OSOTnsouR4Vi
J4bmhPT3ujopdqOY3cYdb8hAM8p/gL0rrFz+VC2YWGaZZy1CCkLf6C5AYUUWPW1z
h+qjQ1Tul1D4Kx5akRgRdOM9ihIZoj6g9arJkDND49Kyc8nIS0R49BnYPiSzdHpQ
/breJhqeVLgl9QeBp/Nh6Xmhs32IjT7e28GaoqpLluFol1BAQW8+tlYYLwTuWIPt
fqt1evY83+HTuSZ2gHy8OfZkQwpsLNGE0lbltj2nj6uQXr08R2+RJ8R1+X5jFOe1
qr4/3K9tzSNo6cIJQmH2//JnQETXKyfgtcU3f/H3UunIqRjRJJncDQ0t8XCrlb/0
LxSRRwmoEUIP5IDt/XGYOv6cZXhQtFpvHLRnqcm9Tyswh6tC1iA8rdgUe+FN4A8J
406APMc/xhHqkec4Hxqdg7hfbPC+N8ZeTjHmGyRXgsxe+LfhnukwQ8yCb4doSAli
ByQFm+zr8jCCBhJ/GXzGrcNFa+AUYe0NTJ20+WdrrWx4tv0OMM6qL3BwtQcEQrdb
T+5/JPny1agqszt0tKB9lbaYmhRtnPWvzAgLaEBo3ydZMtez26qTqwgaXNVmqZhZ
VVtvi3ygfpHVafgWjVrmuPEvPijKa3SPmYb4S6h8nVoqDO0AL8W177o/AmDLkSXy
ru46JwGKaRD1BnpaA7M9AbgCXsHNFt4QUmhIVIwg7ewW1IEtWRJHnDlfNMe1dXl2
0g5biXmbPz9mU+h09b9mRl4hvhKNkiNpRzauW143JtigFOff2i18FPZzs3B79w4h
29VPQNwqHZkmMpeUIWUJTT68a06E7U4jcKd1yOacoG7qsd2UAqQ6fpWoQaiCavlB
IWkEBrQfx5HNz38hbS9dsBGY3k4+eLgM4goE271hchHnwCw9qPiqS9atmeFzg2re
AFXKpyA3txEBcz9aRQog1mQtzYJn9icaMnRAvvfr2s0=
`protect END_PROTECTED
