`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMYUfxKV58xXb/NBRv5TRi4YVkMZAbHJNlgtqUpCpLEt
XIwpJkjorBdTx5rcc79iXyQ+kC/qrEzE1n7wj6l7kg8bwsaEBZlA0lnazVt+A0CS
lDSSdmJzqoYXeoSqpS9prXxAAbwYyKiOT1B0ca5RR/gmaYL54Xhrlzpkvj3CV/ZA
I9H6Hnf1AiiNrJwwbqB0BQ==
`protect END_PROTECTED
