`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
HNESiI+ulhnXqZ+mXLjowP5ZbKktdHnVf+D6pYy+jpr9oZ+7TLTnDHAJjeePqA0k
VBp4XfckOTtfikXo0tY0+QQH+5dDdEUAI6g0LJZBNhr/Bnox96lqWUlv2jq2ZQme
uu6wEt7e+5Z2UCruh7mDY46WRUiMarTU97Ui3zGGAKPaYuCAkz0m4RIV6in3k5da
6eOcf2gboQYf9YJpeexX4vZ9vwSXhgdlD5gpaaJwhcs=
`protect END_PROTECTED
