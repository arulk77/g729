`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJJtVA/SrYTglqNACLkCanch/jRskvIolyWDva3Zxz7Z
m0+kh3t2FV4uTI5pwi6IaXkmrBwCld66S+8eDYjJVCz+JR9J5MnsdnuQp8a8zKYb
CfZDe3EsjqoZeVs/o1fyjKHCpDb7BQKnC3BR/dq1AxjQnwjmo4gnwijbDAtdr/O9
j6M3zY/7G4oZ7yQKSpkx2Q==
`protect END_PROTECTED
