`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHgbdnfXEjcp9Nnz0U8YJONGpoaB1s6AfZ0VO3tyolfo
c23ZdIDzdBAhTzRhSmYFY/M+5o76pXQAoZRKa7QkS88oAYUTUtcbS4C8iS6CGH+A
qjao+khP8EJbllbOjPWWNYMNPBXyR6Qb9jXJLLFgfaBvwIW7xEmCkBsyny+Eq+Kx
wo9eEMcjpMU5UtoYrwMa1A==
`protect END_PROTECTED
