`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePBdaYyIhewes5d9oLQUETXzsh0ZdxJ4zWXiNjacl/QQ
F6EvZk/CECj8rOz2SflqbDo/FAnbLBlb8oRwFh/KgYI1RPoTVBmU0+xp8W3WYT7u
bYVVKo7W+9mJ/SkQraaKo2qVm0/52DSWdl5Zo+9sEkdpFZCwLjjERKAY01JsdKbO
mlHRq04JcJGBBI+J8Y6h7lxCHhkGaLb27xPi2L9I99CG8lujGT7T/HewCoU/MsAq
bsRFNrK878PMYCLJFbgETqcbK2PKUt6Sb+Uudm2j7X0=
`protect END_PROTECTED
