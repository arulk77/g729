`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB0iryY2YbL+o0PUvuGO7dQL1ImPc+jEvl3FEhwE1CVV
4Y9q3IsPPvMWjHi+eU8dVOhr7ykjx9B1Z32BoVAEz2td7K54wJg6BCnhCG6/53Y1
jlK9s4kHhhfFrw0NluZQFm9HrAUXMg2f/VuXV0GLthEdyPsNemU3eQ+QVx02LWqp
mFA2aI3B6kN0xdpUQR/zqA==
`protect END_PROTECTED
