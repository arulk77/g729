`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
I15EiDGkZZbZVBp8hzjOCaWpwhUQ6mCeqyg9ufnNH4JwlacPQhgZbi/Itcaa8U5V
IAWFwfiBnhIs4ur9REve8VD2s77TLlBanuuNEDv//QkDKpIgfKJRisO38GIc9a2h
7JFoqyzUg91EwYvr3Dxrcq20DPRmz+r8UvvXeRK52yBwCIs53WTCfh0dWajCdCtd
YsBwog2puAGT5mpCvS74C9ClH6DMtLAqVCB413slssTiBmYIYpvLoIs1ndTu/9SG
nyvv7zMwiuqlP1H8Zl83dbq4nwtrmfK1kfIWXKTi9XA=
`protect END_PROTECTED
