`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
O5YFUZs/4YO16zNluRz8vAIfJZFvYcnqiM1XvuKh65GOU8upiWL2zMceG2/PAXwC
SVYh9JQq8jqiehICf/grfof6GDfrfK1ip6LmhG/xsdFOnK3scevc/AT7gkXaNM/Y
uMOWbTfQ+HKiY1VFEbikN1peTtqi899Hz7RR70kzdWwpfU8X5cArPsY/rcPw/GCJ
`protect END_PROTECTED
