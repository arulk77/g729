`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4rZff4+HNuzg2Q184WcjftDQ3WKhTN275r/NxvfUrjwwnbJLKird9D1cSe/a0AK2
yVi5lYmJNoK5+Gd/ikGm8h9t1zAHA7p/xywKw6ZOM4mEJoykFu4h0rPwtwCGpcxZ
ZubYR0kHIFE9nUWD7xeDlhcfG/6cQoB6mepnnjcUgJIAJWkuazI4Ulzk58QlSE8u
O3BAEr/z6uiB7hngyVs/di4iAJ3X7JhTJLXnLKQak27DO1k2sfEAohmuP5t5GnRj
quBqFR0aOUEI9lq3etLo5sjJ6AFd5ildw/Cm4mcUPVA=
`protect END_PROTECTED
