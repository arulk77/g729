`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fVOEJ2xaRa35tvkv4pqgW8WYTTpBqzQyvLNSt+ARjrH80UTzC/Z6EDpGP2rRWVgQ
yJZsB8rM/g1nd7fIGoHHNKp8zZNFbc5edGkJFkd12bPstDNf3qBxOnW5JsMIgA81
M86cXVwj+byHESs1R4gegL7dDpqgObLmiAtthXj8Iz4lrw+xllbqxcHf4Zujln0o
vldrWqtWqCYzSOgmFSiH68JOVrE6kw5ts77uCIArzFm5z6tHPmWYAdZIpXM7eciN
rUMrhlf3A1nrjH14WWpNmdYBoFu1ckkJxZqkh70M4jXrxuyG1jL8y3fF/SUH7dG8
jRsNVtqFVnXmzF7PSpJcJa4J+JVh9lFYzYuXeMmBcnPFqKzmXBLTwG8fQ2RWtLQb
MIVUXbFoioR8OvNxAfHBsGeTtQXoz/3O2DmdEydCRBtnsGlHrlUDCAV8zbbimcdp
tzYXeq1TN05bOruRpZn61oWJfnhNOuZUyZ0FQDX7YAY=
`protect END_PROTECTED
