`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ymakm5NjQNeTNEAJyOvjA60BNfHDUJKu10+B/ZVC+3c
C711DJoBSpw+/QjPRmw9iCZ8mXJr+p26JrCoRYaqB/ZwZpY3XCUfxPrjlJwlE6md
PD9hrUZgWjLBO4A+wbQkhpxycRIutWrYaGiV2gx/2KQfmPMJupiHJJCu0jbTq/8+
ja4vcpTNajyLHS9eGQyQIMmPnv4JFcNCZf0r01Y3Tq3pU6dBkjrcRCSz3oU2AAXu
7sN75UVLa8x7eYWIPJQzmWTQVYsxqnQ9vCrokseA/L+kWcgTMZPdTSbJjbcUBH7O
J/U9F/gHCims2554mS1SQP+3s53lCSxDiYGhdau5+B9E/lTLqGodSUcRzhAWPcVU
t+J0r+hlZzALjcvwTeDmmg==
`protect END_PROTECTED
