`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48kmA9rTXS7w4I4rXEzSFu0DGu0MH4jIgqduXVJMCuu6
UrTQZqaLi+TvwMyqj4qgRF1eXWb9UtoW1A8Tl/HDqfxmhK4JyRxITTaDhcgPrHuu
QGmr2W09uuOrf6bvI9N52IVBx7bS2RVrCUlcLwadtvMK8unprWAB1SKeJcOdDEKC
hHr+8qJy+mFHh0JbevSGNAQDw+LRmcaqgGqjWa5Z7XVUpx3YNU8J4RC1wwatXv9W
Y0H5z2tGCn8f1FCLx7YxejNZtAwQwXuC0bwAoO6GWbo=
`protect END_PROTECTED
