`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SZblvb1a7RAY1wCCKTuTOKkDah6D4I7ABh4VqaoqdjrM
DGx7AG9UeyaicZU9AyazG0gMSYx8BmTZObpFk1OVhC9V3WZanDklADtzXkc/Ou9f
x8optBiTnb4y+ksbsCSojEvBh4ta/6XHgz3Lrt+SQi98Ofz1fMVcqNFs8JP/FcVz
m2baTBir9MJZ0Teqn9Yn/w5h6UJvU90nAShQ+9dNxfFUR7wHQH3mT0DM5SCuirhH
gLrVGnN+kwGRZqVOI2oX3Hf7OgNfP4nanEKC4rsQnFKZDZJrTi/N7CgKWqg4MANl
q/baVZJk0lQOOThYNIltC9zvoQUK8qTrGFWJGc3+z6SBbMF/yAlXCtyu2QLYrfz+
+XBuhQklclgsXwqQDBqWH7/8aGoSJeATX0N+zYctk+ZrjxHiqUZr5GA/DkOSofMB
De1nJYjOpD4IM/rWTabaT9+pQq/zKejYLbsvW+Ozn1igYqHmGi6FWmuVsPv6lt01
h11Y3AiK6JCrjDE/w8xMhlY5iQVhAbofVNQhuZywlCLTn56G0aOe8Gsqge0dEt2z
vJtuCtSyy82WHmWRdcE3SHfpauPPGbbuSVEqVRm+0+Fsq9SZDvJa0dwkaSwc7AH3
k8ymN61fL7zTomqoD0kojLR5yURpE7Mo8rglwUtLuWQ+OPct4+i7SXLo0ZAdYswW
GdLsDoLstnyntNxrmivrD6NwLcgxtajOv4Om701SIb/8/qei7YiIH39vfJGsK1Cn
EWz/hDcKX/1IGRRUCIAGcvVghVgCfCbrQRzyJ1Hf2qsA0A2ZZIh6EqZ3fUTrG5Ds
trlpumqdi2ygQHTk038gXGliIAwtjbfrColwPGBM+LswyL2dtMYK1SKg6tTUnqAc
Wlj4nSUGCuEOujL7jGeXf3M8irN6D/IpzRIuWIN+qUDzZHT4qDpTVgxTLcnPi4m6
FOxbsMM2L2oM0MoEMPK2CbHCzPPbGz8Rq4Ekvr0yuL8utRc2wTnJQ1w+2yULUobM
z0ZUCnIVf8r75+HpurlA6+zcVLUBATV/IY05HMqI2WQ98zTtN8FhfbjtdRWpnksF
eZT5UhDMm/xCZDC+plP56p6tBP1KbqgMKjZylDr1LbCT6sTlp7Ms316ZI+zsvSg8
Wyz6MT7XMzCiqSIQAXsGA+9ZV0Mf59r2oL7hpAk7AEg0oLNHW8WzuozulvJKnGn1
PbheFdHDa6WMMrZGrlPNtXYvk2lvi4QO3Yb335VLlE9gQbHgxm286kqUgMQpKj8V
ttWfplL/EQWNXcrRxsg85svbH0+6q4oLKkg5QrVXuIpiaXym2PolV/32k6lnHR6g
L5gjMogUpuZ/+OdzDSfNGJ0XEOMhdHSBJKPwqaSHlwUj5rvuIdrnbfRio5jWecei
ltleRuvCLE/I9X175tZQFsKBMedAkNC/kmyTMmzYsjcAzkPdC4FO5JWyLwVOcBg6
UYOtNZLHcoSOa4oRu37CDp+IsMVdZ5Hjy/Qi9gbJe3EOG53yZntaHr+MRZDPj7lP
YYpymLR29WmWXscc5B9B6rvFYjuLLMgqI6NMChhPFUDsDPJEYIHmfdFBaXUPk0zj
XMn7OqkRxG5mVyjZLSWGbywWX1++I4Cc/afcGS2lb/vGO5hznVyHUTLUsN/14okD
nePxVDIQHVXnMRv3m3BIFhapg+DY0EeBlO6oNSZwXMef0nQ8df6q49Vc+URh15Yl
L7eXdIqWixfj/ryeioEk3Si1WJ6GIN+MDQGRw3D0SO8XLhvyD0WqjBdTHruNPlgF
cNkjXE25J1Y8RqG1bluVn79f4EFQ+So5oel4bhugDGPUYbcfvfuPQJy3XmQHOOVE
ja/Lw4gDyKKfvFuLMxp8Kio4S7amfv+YL9aKf0v66AAwKSBFvTqVH8E3j5qDOnjD
fGX421GxrCQSK50cZWle+AuZLst2u3IZwjk/hk6mB61lbRaYTWwNKfrGFUaWJMxI
+UPNPlpMgydE/SBgghXZb9LXlg6CpGXRwabHy4OZpiZQn0RrRktMHaXWsAK9ULNv
z2aeYnh7LqN3U0OSJnFHcliv/RiomeYICttoq57P9VQNVaxq4vg1CdEC0sSuZI6V
3yIy6rc2/0Dx1J78BNTvtBFL9/3KZLLE/+hz6B35lvEg7X8j7pDk2NZiU5o0hHHg
2muMx8uDtdXzV1eti8TJldm7QrvC/82msyHL4Q50AuaSoTt4XfEsEE8IQaCJLCUw
RUYJ2FLNKCzpzX5BGelrQrlsCCvnWQo7WQ34DSXLJaI+U0YfC5wVobIqDpUh4Ith
Iq8w8PNc8F8HURHIFPNxkuRDvgEoHSs9GXzw10HLhnU5SWyV7A+z7UWixSfkGJGG
8hTCQuGuVj8tP/JibJtJyVHLjIst1Q57gRBTu5lozVD2eszWS6ji755rAioS2RZa
Xk+5SrQQqGuF/ZAVakQ7XxAZl/s92tONX3taFKH9EL6MCQPRUp5vjEEoFSrCMG+v
lBsdpC7N4SarwWZ3+eQgMmo/m268nFSUQJi5PeNYSwydiISbzAH7cTzBcfBx1SAX
qU3smX2AITajnj946Z1v4bRVKNPcob9d8dXGnyrO2Fa45OyIYQkkBSQXa7TU//8V
W60uBq3JwI+NQITbYlOG0HZPZsTejwIRH9QnbDsAiLLeSIHLbxklAClfWTxb96jT
aRBdvIUTSc7fCF4/Q2ERNxrE6wB9VlCUsD6ey8MUJP3SscOLdpUfMC8XpF+QqqdF
0RT+9CRaRUtmpvx78u/o05EM9SSTDid5rwc0NSi6GXs55pNpGL9srZfUphpBttaQ
IVvSn8gh33u2mFsOg9AK87wqc82675FgKcOXDzv6EsaEPDn2PsZ8yzs0PLH6a1Sv
nuNQQ4HL3qAXHdX5up8aAGMau3SCy//AbXABJgFNwQXjw14I25rhC1nZCIF/4q2E
AtjFtyTQ2cUpZ5yHGo+AarI3Fh5WBs2u52wgVkuhbD/jmAAL2tcv3ZMJRi/3IrHS
OmS/wZJLJkNoQcMKgLJZex2H1kWc4zWMewVAxO8zs10DrFu7YXSKHfTDma2g6FCi
w4DSCTTnLMWlM53vgN8jQdPqMpeLKG/GIOgPbCVYIH+HC5tNNPhDxfse3sl7XkkU
1cE77jCsTkiS21rMNi44szsqbrXckvIbGlSZvkv3Uqduvva9P/z7hl7ptQJYeE6e
zgkXRntNMJFUPdoEnErhtjfrF2gO7RL9HOQwNCdHP53AQKIZ8NWO2N79Pru3PP0+
6rjbcAMW32q5brjuHA6TQeEkCDOYbjpA9L/7hkTX2zeibKg2acKX1fY27KGNvdEx
zJSGh4tUBNl/KyUZkBrSK5rZH96fllI80M/nfqD3DFxQaKQ0Qvci2uTlr29kjMQs
0R1bye5a1Peitfx4uPyyMg/3n9ct9PsSEzrciTqE+aAMdPMTawAW1ewd9Y9TEyk+
nLRQSJI2Bgn6cT9fgyIDXxsFjbQNYWE1wVO0qdQg+JOM+uyz53KTs8loTcUi5IgL
tqukMzy6VgdtWxclR6RJk1neapBYFY/s6SDQTLT5olcLcExjhPA4Xe6+gukQn/bv
MRqmicGrAl6MJhIKTYiXZQeWBj77ECNS0UqOKj0HIKNWDJKXXcpFG4n1gefI9rRT
2B+B7FBEEqUNvRg2vaT0OjV++pvG5RLbST3ixjmKyu0CBUIQ7Gsx3lHFijs26XzE
tRRgPfS1jPLxJApRdHhu1jDvbG0KtAaTSFYfSxe8QWKRONUQVEpCf48p5dmDQyZo
6gy/fy3ERzj4SWyBShzlASOuy5sbHBaB7SZ/JNDVUlPV9oNo63Ny9/a9j923MoWw
6tb4v/NBcHWnmniP1VLt5B9VL8AfHP7J7g2/r4tJSWg1klk6NZ8GMw9q2XN/+xEv
cB9r6nnt0l3eq0YjBJy+nWxS4zf01IBGIgYF5QnukG8BTTk2BhYLVTv/zkuT5g/V
QJraRJYPpdPen1XgPEK5mdR+QZRgFurSV90RiYMKdYdNWLelSwN2p5Kh9jAejWMQ
0RnhlsP1VDVOI1zXdI6/8OTBVqBqXW6Kv1zhMj7LXhaMJ5GlSsOjrPh92WmRJv6Q
rWXvui9MQNfMew3/jFnmZ7pav9j5snHGIqfRfL2gagvC2RAMVwQmxXoOMLK8PIIs
x52pp7z+TS6Gj3bbw+oMiCb4RVD/NBwgPmE2yoRuJotMdi47GVS6iCtBtceRp4Lp
wlEJUVAtT3Y3wM/Ud8ElkvmGsDqXnZcgWFRmStH46SXoui5oCxLVaTLmXkvw/VSX
3ciL6LUV9yVqcoQhmVbxjV6MiQ0WU/1oysPwTSgXbOiaRzyaXHCZujT62yCQkJ6E
tIr0T1yFIK7BCEvhl3f2U5tAsOcXqoPMNdRMcnDlVgchG+Thwgz9ltnlhtAgsTqG
doszF3C+Z+8YY92fSLtxyqP58ZMF8ojXKHKyiENvPSgYMbezrNQXVU/F1J4ZxYEh
ANdYV6U6ndcuMX9kamz/k3aNatehvdR6epfoF5Tt3rSMSPIiGEsA6zFMGajsi5ty
5+tfCd/K7o7eo1LkT0n/FuavvKLtDQr5AQ7LJ2thjNm1t2xv0pVTJMq8/D8ZMZZ2
cRy+m3LSQSSyIHxgvALW3UNong5iEMAUNL3gLRk/0taIVzKWDlx2xqgKdGwiU0v6
pueOuroNyg2KfC9FU87DKz6XS2kIhzdxpAsBjUPIKaQsLDL3FnAjiypQ1pq0ydAn
l6u7NCjXORR0OCSDzEYTfnIZL4dGfZWShduhz3apzHDrU9CuefujIxlkQj4amFpW
1DBkoIoCK7U+h8iyLrjulZIzUgTjgsIt0tRJkG4Kcv/qiK4AZ5yiwcLEUfql5U/i
UlCpI/dpyiVo+r8ASvSIvKdTs7K6z/plrn9p02nAve73NauxpfyZXCubIoktOf7m
qPjsnsyPIDzBUB8XtgMdobWiiPQmemgwGeiH0X4N894Zh+POQsbnegM9LUnH6FVy
hv5PVmTt2gpMR1+mQP1BFma38N7JZJta6GOyEfToPeRxb1KsIjkp5lSTq0DlnFtW
hfXowgeuzoNzWyjNyw7WRwgyNR1Grrz4b9tNbU4kv64qQ5LsS7U4wxdnTUKDaZ0O
kO6u4+6TaHFgeZdbsCmhL5l6bGbGaGInaGwZors12wIVtptjt8i0B1mJhPRroAOT
DQMcnwGZ1JdwJrjYBdnf085fn9iuGDkddBshD2tDCZsCbeizEQIglcWPG1oqFtpO
mXOC1jaZXN3BhsWktYms8wisOCWIXrfI5wjH9QN0tBYEsPyI8UK/Mnewol0O2MHK
HNB/HLt73lUjHfjl/DvvknhHYLivX72Xeplp1f9Q0B2Amzcz6I9tGZ3a3qFXlV8g
/Q9u2mhICfwp7/lT3QRMLRKi0Qi/Kf5wHFxh3IndNoFqS3iM04Q6/A0ghF0E42Mc
oR9PmkfFkPdH5eepMbE7qOCsWF2+nz+xw9c3vboB9EAqGlSwNFMwjyq1yeMy+Qnh
Pyud7Q+GgdAAXXmAOSHWO1iOKBz+H6AGyLlLUwpE1rXtbsub2o5gerUaRBUelEW1
TxE/UUPM5IvsZl1sUL/mrTPJ1udd/PYytZmdVdL9I3GS3amXLTPgPFS/lJw8r1UB
3h0RRDOAm91MDXtMah7HPvv92UqLlrBjoI8Fen2rPMsUjDa1lPBFr0AYWDeWhMg2
wqy5VN3NLyQukXAFNoG0/eNPk6W2kMexv8aSAkC2KG3+JARmQ1GybtTgFliCasjI
PSSgE2qG1IOiNKBoblWJE9Hg/x3i22iV3NHBhUT5OyXOqKVNEHp34T1nhbzHe2Hl
tMvwqnLWJjtVP4aP4KO4I0KMv+gExSbSzO9wOdwja+tcleRXYm00HGNotxAW58Op
aP8hn+n99SBaI4GGKTxdwDnn8cvzJgrsPL+mo51Z50p9WePkiJqVKoe+acbPd/rG
0sI44haD4igiQtgvr4TObu64hjB8E1BgmAWqN6bAycNqw0anaZSA/QSq/fO8fwks
AWlLlEs+RC5eLwuWlwpztf4aI5jhXGasZyVis+hAEeKvdxiEnno9kw9eGV7nc/nu
DNp+IkZuZJdXheNrOGJjJi6FxDSCOtLL/Ileix1bGmPq1cF5wDCGnMhN+PIX+CSE
S14t6xEfA7BWklizDkcj35/N30VNgh8Nj6haTXIAK0kgXFHYI0Gvv8rbsXBiYH64
5ulCbrQXTUyn/TwSxEuhEAixcsIrhTsklPgA7zBnMb7dG6yZpsjoS/6nLklgMPmF
DxDUmL2iAaMqWkcGa2QpQpbd1ZDA/z/AQA1glrvtKBgT3+qy6s0MfoMJ8p0B5W2p
4XlV+7H+W1dyMLYgDZPc9xvdYOKSvy5RfUJtnYWZu2wiJdulhJ7k7x9VZgrlo5aY
TScVuiiw7j8d9T+9xZfiOmUSWtXtwCdC3GYXX8W7hHAekIziqlRTFkAWU/3ftl11
rT4yROA2QRSHyxJq5DaJ+YnPnRfCvNWb0ZTdtuuVO4fVecU2R+GzDxJRora2wyi3
WD7qOzg4upkVXTT7ikznJ/S0L0bXOIVXQtCbmherhaMD2gCgg5+UmlNCR9wlI8mR
cq9d+05VJbJMx42wiVmS4SLEZwDwgvjrbhFHCLq5vhs=
`protect END_PROTECTED
