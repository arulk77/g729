`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SQWx7RZVPaiI29eNFnEvuwtiS5qYvJciC4F9dXNetkkO
LTpDzWaaurSFuUNs6J2zi/SZs9w8WFtgvyXoijtkob21OUtM/AbWNmYdjhZSJqAS
/b+GSTLV+b53NqC1aF/mtkWkJ7YKB/SzaBn351fLuLbY5CNnZfo3QGj3OFFlBkf9
S5/rDhIx7+kQxwOJaP1RVLPINTpNNToxkTDO+IHajyML5Q6EDlDuTaQ5fibA0A9i
DGdcgbsaiSw5xBlBH7F4Q4IhXycv7osoS40rX6qL4vk5bT8+soXFusy2dgwvVoZ6
34ySRH+Sgdnb6XUiE4wNbZCu+NgugCBq7AgI9bmYVeClxFzb0tRvZNipZ6jh6sZ1
2EC4KI0JbjUmzE33gUPOHjQgrOMrByb91Q94sO+87NhtXlCc71x1J4/BZ6QEBiKh
TciZItO9LHLmqdQV26JyQRGp0rzW25bk4dvUQQOaOkkYtdRx/sYB2a9FliJZJHXF
qo9x3wU4N/ju6I4m+KoWkocs+q+oLenkAgeqyuhC/VddiRjX63XI9kf5gaIhPKka
LdCzg5dFAmepch08c14mB7oj1f46GH8V3YOCQvTa434cg88+H9gBgpbngNgN+EZK
scjX5cE4bg6hcPkVmN5x2iAFlwpKUQtpzNhE+LzMzkHNA+AjownfdkgLaz1rr+pz
taxrX62KlK3CU5jLjWDE4kVWBlvROMYf9FqObRUIgO5oyWC2XyhTFvZ07aYpmt5K
UH7dLsNZWwQSFLo6lXJKBuQ4YXCuXkjMO1WGQwbL2xoTfwqjBrWQZ1wSgjKnAmtW
WGktaRwu3BARVT+i1b28QuXQA3T6u39hc40VDmDPpHOFf01N4SfN4v3g21ApLFWU
KFiksvNvOFopH/AepU4ElGFhI+EUdCPZA4E8/cLDWn5b9QiTT7K4yPoReLy0GNtH
CtNstJ25HRgJNBxur5c8FezAv+ettio4pM7P/iZWxFxlkAW8k3ZvdxXtYxYSKnbe
CkLR+wlDmjyrLVxxZR8BeqVYjNnZoIDaDJLyY3NhqmhSdAFYmlaDQGn9AEpQe929
SpnYdbDPpsz1jzIaxDjsi2YdxnqL8JxbL3U/j17NhRddIqR30CeEMDhjvnjcYvIu
LcaApKKlzpZ6LwZIHt77hCXj56AjiUFysL+2Fciztl7w5SlS9EBRlYkFMboE3ntJ
eg2VQxBz3zCx6MIsRLWnvQgKVcnLvmyVvz+tG8oSwwKWW2UMwEtfajtI1FMmoMSj
qZpXernfHixEDzeQFITw96lXi5c6s2A+3/ZbUecSUogqFQ0tJMyx4rKaPsu4BDnX
S3gf17si+lYmfVeFB8IexZasQiadJXvvejOCc2lTRhUdkPg5mTM9jFzWhLrNuU/P
pEiIL/HXNkdnuVf1VVtTTvCR1968ZlKlZrBIu8aUf7KX3v2oXgVZwGnkpEeHGzjk
SsssLwBQDg7Q8seyDWOjdlcS4IWL5dDSl8qlQ4ZJKWK2XNLY70RXvLjXmqmY7ntP
vYzWim9cipHyYF06waj5Rt/6cNzzDeNL5R4YHIcjlSS6TsnGjpIdaT/Und8yglbI
L4FFNIqv0CwLtN5GSgqwZGtwIxsteyqL9u0nQ04JeUDuvP3x9Rn5CYI2MrgSYkyJ
Sr86m+UJhRKRWbtrOSGb9hNxOWFNXvkmciZVk7iML44JGl8fdSQuAikgHBtyqRVQ
wzHpc2ukMjVfkt/JiuyD1T56Q41fwIvoCSCtVs7JRDlWWf9phSHHNE/IP4rcF9Yh
IMBruFF7dvaPSpTmByd15b1+bKD4bDr5ZsZ0tEKhYJy4nvl2u9ROV5kbNsT8kXEF
TBxedkljj9my5ijR1YWegSeDqCfJ3me/6FEEHkGDB1ZLhgT/BROtEO68YJWGg8c6
L2ERqJVZV7fPsB8ZY7psff2BnSXySpUIf74GN1FYNrRDm1n+PhtcjAkxDs5uy6uW
9gL/oXo16E8lMkxjRWS9MuUBP9JG7gcAlsCDa7tOEW7W8sRTh40cO01/9J1p0ijK
5VrlT0zejxp/sq6FD+LKc8RRDPTfFb7QfCbYtyr0jnLW/aPjRbM9PHOEiQQaVZBL
tEsfuDO1OqvSeb8C3DGSmd1DJLbcxWpPcR6YpDpIIRSICfUD2c6UhBUAaPsjInk4
ROIYRunpAKkt3gr+nXJFc+S4BsEf8+Ia8JtzX5oyaIxVHQ2UZ1VhPxrz2y1WIDkm
EQ+O3aQXJPiwFrkV6VZr4USlxghxZPqqLPFC96xuuk1/G4Ruil0jclpgJhsjlYrL
i9davx1wlf4NSQU5q+FiutN8D54cU/ZmM29X7as1FYnPH3hGg4M58ADOrtJkklHe
C61u/iuqacZVVLhS316t2UBYNfkat2PS74C6JuUBiTBkW47x9xofNkox9EvN5qvg
oAuI5R1n/goRbeciVS7EP4twxgYKD5GH4NUNuIA49+vuVXayY5WdxJaolbLLZ5Vu
dxsJCcLuaD93Lu55zUJuFBUo40AOtTL7Zf8VTCYsI6KwE17yMTVWwVF7L7t86kzX
yL/dqXwENw76VO8UiEfXy1YGUnUojbST7Wo31BsVtavgmT7/u1ADf2nXQ6HXXwCN
+mTjA/vtvHpuPumintKmSacKSpIVpk+3p8xlJhZVtFYikYTEa/OjGY9uIs7F3D3D
Eq2PKzT+w3o3HCGfqSPtpNtjvjYT5+OEdDoHAhrrUmCDje6qlbSu2fBN/O4sgZPF
Xq593ozRR+HxI++fS6IrGLlP4pH4po8YhUrIKQA9CUl8JmrxcFJE6yNqmhHdoBKj
ZSm4Ojpk8RwMVJuy8znILrAKJVcSnII4I+3P0OpZb6sxEsOkjiVdvlK8+mTizuss
kGRSP++chr087m1S+WHRUickv+ihE+zz+6px8ucWJ+ZBWxqUzRQWvHZQeLbmvGjb
Enr3DM39TfI3mLqJhc/k04N9f5KlznQIezcv+LI93QPhKYlnIosaZeEsuiMF1O/k
+e4iykRdvINO4k9dEMNI80Q8H04oGAf1vqbNrfCqE6nPN5myetcrDTeli+2+h6h1
XqGGCl+8pUlCUeYJxz9fPCvUPFKDjLeB2ND/1rY2imJVJr5TVpcST5IigURo/Ndm
iKrBPKpZRNfxLvRDDAF69WCx0EslAUUZQ890ID3IGAa9deIB4qEWUlcU0O39OQfw
z/zCAIT9BHQovpGnpH0nPR6j4zFmh/XiLbpc2IFK2ihaSStsDx3lg72Hx/7ybxnb
p4wRnQv+WAGmh+6H3wdCendVDi3/SYSwzoTqPE1Yg085OjDmy8wGekYFaUY6sZA4
51FDqtDmzDHfd+tiiQTRq168b8q/ktiX53VXNRaURN571YfXRFDlnwbb1mLMj4OD
6AvUFPTmhmEyOaGufQndixOqSAK5STd1mgQBkjF3dF3SOlgr+WF1yCqKJ6bkx0JN
NyAhvp3uqxEjG/GtC3lcFKYAWXnck/htr0HWgxz39lqGGC/vCMA8PEMjARjipO91
+WkbWovAwJ7cWQrAG2dfVWMn32/31GEps/9zPnTg/c025pGm8LGQ1mIyEyfX+/dO
PqzOdtONWXtLId3x4/clCMEQUBdKFX9VqgLS2wkb3IV9ObCWJ4EhTLFRpxCFb6nT
OuOesxR5TMwRTRMYqrm3bAGoD8EloSwhuyZg1RVUTc0E83G5ApdFvzho4CsdA+1t
8xr9UYc1WY6xDjsRlEHSYJ2fwGN07k8Yf13S2ldAJsEgoHdaIkEKD/45i00yNBV4
qjs5OIODn4nshcTXFeokaFvMr2Clipmev57TTZVClevdkBq3j3dLr+b6qWJ1glfO
pSVfyD9EVOyUmca9IO5Hr1vjt34l+VuzqaY6GM/KYD0KmPJCx6xZmX660HOaSBu5
v8CoEZVOA3yoHpsFM/7eX7QiAgkAYJAddabz8Ur5GaivboRC8hwgAyV5l5rcyUEU
NjNaNxuQegYgd+xLpIsJBlyPVOI1LHWH5q2Z67LLA2alStingxJfom8jTqLM9FYS
THiGrWr4mno6RU3Arv+5UsWNv478fzQj4hikH6DwALmbXGXDxRhopGPcOcWiiJPB
Jea7bEZgKQNpMvnnCUIeFW6YJQyDG5ASqKMnfj6kew/e8/uCkhCUB2ymwZl9KDaG
WhcTg4vWh8vH9Uhxds9mZpxR6o7Ixo3yTQdo9pWHdetoNixWpeD5QX2PIfpkiRql
J9nmFOIlJpjOOm5A5jCJPwganT2J/yrWBPffj6WJesjwoKQnqYk+aF8z8L+XaV5e
fYJMX8XkQQSV0yPSEQMxsUaeVEwdZTqMjUfGSWQqk1Ie66F2nHJPme5YedJg8SX2
MRfLJucFkdCBu1KjWFEzifsv5lnDPua7h/iauWmNkkCvePpkLulqJv0xUARFo5mm
MBkiwRqb3LXuU4Wj55l50keJcSo/Tb9gGwg4km8b2+nSJfp2c/K6lfV/9qbOsT8w
tYp/mwYyOtJcWGPCoEciagLspfQwbCmbjH04X9jg5a42JJhIUoy27O+U0BJUQOLS
zz5ZwiTDN/NqfobINDkrvnpYM+99E+0CrF8xpqEFF9E+0BhHm+DuRNFUfkapvThU
inFa1VLoV4ABbk0n7ikvwZqEbtNvnA09BeSJC3v5DODxOJPg27MPhWpS0w6+TuR2
cYw32lm6xAISDPKGhtY1W1f+EFIo86ejHGLn0/LZOv+PGkQjutiba0t7Lh0Fl0ph
O3ki2YLyxXF7aUcMJNyLTKEnVtaF9fpS9J9DBcQ0MohOvSB/sFEFD3QoqA0BrKsB
OYFBIgLSFf8jBz00T/8yNwoMeY550aG4ds2OnQXQTjcy9ALVBlxkN3SKIwm1Zv4z
v8SUU6Y5HevlpiYUcncWDsIrPI4Fy4WLNJacdtMbf+E0dRv47axeq+yNuob2M03o
6LRTHoecoIHdxVGYKdG9lLCwOuJuPhhwJT1TGk7Z4pkmwrs4c3TrXVz/G8ApZWUq
nzim9KW/+631SsNH1N+Q1F/bwRWnOQaRLUQ7dxS5QpxMvLG89uxtgoBFTMsB+iVj
csUYOCcpuoh4B0e48Q1QIpxA6LCBk0M43drEiskGDiraExpSDEd+a1L/ybsgfGyI
6RFCo1pkqqq6bPm9IF40DSwjz8NNkkxqjH0qwt3AhrI=
`protect END_PROTECTED
