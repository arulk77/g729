`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RrzH0jTUFVKKTYC6J+DZAyvipIDKGHQhLwCLI4tNqMDl7rTM8HcHtR1dZ90PP+a8
0XDakKZClQYfVOk50dB6vkn0m2x+lusw69A+Aqi5DVxWrL27dJBWAmzsLehnsQI3
QDYKRR7jKiz06Vry/Hg96Zq6nTuJdEvHndBALPH/MTfXAhdBODEwwRsF4RBFVkeb
h40IK/a5SV9jGvkUsUJaAR9hPMGDq3o3rH8XTn7ZDdd8+CovTn3T/56374QRSpzo
HfW57QdEQgolDirAqOD32e7BBykM8NtD42YrXVS2AZH2PxqCFwT7emWSodoEVjvy
1KLo/zoeWLvUcAgmq+GwFf64+RpQNlGcYoElgMtcXElwYyEU+J8TpQqfcgoKVXNZ
ZTTFEBzOTHTPwzVhohWgpmK8UuyFHDLug0L1rqGWx+U=
`protect END_PROTECTED
