`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CXDo269tkFVLssJhCUcbkZeVX/pWI4XGhH5wHvgxmLAgUWaSEkut+e7B2tQ9WwiX
D97LYLHSWuQaqDZbQndUy+YMqMjtbEdZEP0o9lcZ2hBM/iJAqOOInctUd+cwH5w4
PfaRzkjf+mB7YAjDTV2/XT71YrSpjZCbSSZez2Bi6XjCotUbWRQQYrg2b7S0pKXB
`protect END_PROTECTED
