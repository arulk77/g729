`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ8fEAulN4bwDCjd6kXT8aSxU12GPBbOVQ91F7Q2EY7T
SnESmndxmR0NFZLprvT1qiYradRvevVhcUGh6KiVc7vuDEE3acwj9DuZBgI8DxaG
a6ya4J7/tOg1ytGXDzkPiGf6AIUmld7WJjUEIwyW2L04QFw5vlStqdOEckLxFci7
itES/FZveRgcCayO5Xn7xlLyFVl9bREv6FqMTK0bDVE3BldO5oMKmzoIH+gMkJds
`protect END_PROTECTED
