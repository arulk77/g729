`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLi8ER0i7bONSP3QBHuj3bk8wgkAExbbkDSPbPSI1D0x
97eIEbBlDu0EerHSVu8G2r2PZlOkeChmEy8mHGKllQ77f8+j3xsdCGFXS/VNUFLC
cZFcfr/RT+Xm9Yc/B8yqsfUad0TJs7Q7FewZ8U38Oivc3ziKXBB7kT2Kwt+1/Zbc
+nBHicuhEWBxWipXIeFWsbaWtRdB1ftmWIyc4RAsfv6QHIHw8hiNT6r3UYpUf0UF
TwnnZwpzrPtvCQPYZAwcsAgEwbqGKp42h4V7p2ouPbFCYnuJqKeBKBuoj04gpBFG
4FDi10R48dCu2p4A2aRRCCF8kJg+PTNptt1k0QWDpqdpvZBWmKKMxZ9M2iEy7PLd
zpuhpOqf+DI/qP43EMg3/wDNPuj/DC5BJfMIDa4iqG1uC0+yiQ81rD3l+Ut1zhoD
RfDAUqypF5t/akuZ7vFnHyTRuTIl+2uiKZ9yCgDszo8HB+Rb+Ry4o7pMAEcaiBeq
TxdPrC3cFiVYMU/XQqdSKSh7N4+V/L3RVhPTjlxxVS+uYiB/LgKX8EyQQvzpjBSI
ckBVg6iDFn4XVcwv+QEJ1w==
`protect END_PROTECTED
