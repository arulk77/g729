`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48dket+l+1rD+mw0HXfvj3dSOOUPXS95IKsaSwE6Om7i
VuCykzfJ5Iu4EaSpje3ZrfjGTjWYSCs30e0a6xMvOmVoTe1SLgVwAa7CHnGaD0Sq
RYL99r4D2OHXInQul1jQxA6+mbRoqjNaWgRceJwFeRnZYm5O9UHvQzSQKpw0afr+
2zNi3a8aXXThid/wZfArbxDkqYdrWGFuV19Ysme0AF1CmYhqZ1Ith3IL/ArzKIok
lyCTO7wKu/2nmlXY49+X1vso5o/Nc0PHkcQlNq0ndAfD+KapR9toyUFhHlzUYrb3
ZIwskWLCeP2MNxlEeaEfQelE3deOZ4DqbF5vCmsa5FEHxaUj1XBfBLxFdsunTVbk
lfKWOZRAUUXb5vspOnOxzdn0XkPNsrOWCGnwItbYzpakAmQrJ2MBcg7USfSkdimk
dHLrh92FLwX2e2GcU4E8ymUBMX8IfRXR026qL5EIXyTekTj55Ex6k0RebeGSqaJN
iZabuxflfrDY2zdT4rzqbPsdwIxgbgrm6D5DyToVxqxmEIY30Ip8aRlbp34PCK67
+Ljf6xR/zMmXAT0XBSwMClBdgwEw34YhUsc0YSdYD3ar+zaBe7b8NnqkbfDNF4f0
pP+u9PD3XFb08debfNva46ochkQXsz3b0AMxUWXsJO2nf/Hd8K69p72SqQfrW5XK
O80hISoJoHnID5i0PyIuN9jtDehUbea3QaHm7i1s16X85TNpvzXNgUVdXvsr/Bjx
KWZ/WG9zCJ+MKKYVe7fO7/K3H/0sMdQstdBV3PefVuJYDDAGCR8aQgQa8RX+usRR
Nb1oMw/6KyEt4tefIjmxYbo8o2O6UWHPwZ0RaVb40q79G8/qItFUEW7+apg9TXPN
HVv85QTtKWBkj0sJc3wglm21zXkY4ZMK6pUnG07kdw+6JRI5scT9NfTY3nlB0Oqr
/Mk+r5ZaJyK/zAneU9sSt6noq0IEHQmkSFK9ZWmXj2Zs34wVIOkpHaqsRLAtohKq
J7uc9vDfxPk4ZXCieZUWSUpvTgmgkVaiHZ98MrxKGXeUNsVboK8QHpM8OeTCSShG
ZOuPxsjUdixm1wUSkHbhDWPPqQ9DWdwk+cL43fBOeeDW44CeKC/g9SoZ0/lZ5C7F
/GlnDB3HXhPGafKIyt3Nak6qid7yxH5xcjVb6ZLWgvEoxQzGzrrw/OL0R9F/OVVs
cU6nPQBah0n/lv0PaNe9zK1khFUbIvie352uJtuarlArICkd6DC2CY6xrPL37lF6
WymTpKWYzUKWLeJh7Dd3yJwUeC6GmHT6BmxZXA16fhg=
`protect END_PROTECTED
