`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDa4fmiOB9zfQ9lLzscQ1u8/UIkBkuaYtCmPWXf2CURL
cDiD9RJ8R/IVwiItqfD4fxKTBnfTSpv0/VZsf3/+nw3rC6AYw258/OoQx4DVFX9Q
pWIB2raq8YEiEW+uewFHdbSoEI9HrXiqm3Q88JVtTkwWacGXqx6B3ECGkm00F6g3
GXtsDFPk06EmO1QUNR9y8MzQnWvOHUedDVn/zqz/lPOuZrLF9SqmU25VFi8ofmBe
ppFKEwahTDUVinJ+AuRQbe7f0Qnd/5OmLv1tmJP0gS6NtdAQ9OmRH3v0ktzV85n6
6X9POxWlc8RLQ/0jzJinlG4A8/w9a1WVxCcGU5YeWcN3mb4Tio08cN9IS8lpQ9H8
`protect END_PROTECTED
