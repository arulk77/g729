`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAfrcGbOCv88QvAkdRRrb4ApE55P266OQkLaZGfMBnn6Y
r5XzuQPP65GWhRV75Hxgx2heR+YoJxv14REhJWW/Ws0uB8Px7YWFmPDGikBblvEy
Nza+dJQtB/IWBnvCXynhJPrUeRxL5NmkGEmH3JBEsR3fBPIs9YO8omm5PfM5+PH2
I6PJdlsz6AxvPGkUh88OrowehOVEpbeRzQwCovygMGGllllXVydmmgUdfdmDD/Y7
nu5k6LWZztrGyT+D9OUSmx8Aa9JdoUnhYH80Lv/M+vonzVK4Tqd1NDc5b+oa1QG6
h0JyeQ9od8W6BCoNUrEJRx7rQ5O+FjazktmlXIvE3w5yJ1z0E4yHqbbATTJdpym0
f9kjcIi9L5Vqwgp7d07HE4GbxBG4XeP3j6WL0/e+h/rymq9xZf0JUTw6BorHhD0R
lChJn1gHN+ScieIWA/0d/MjV4OjPqMRBdfGTAfORyBqY94LEr6EU/hFEIxsaUSrB
AlObhAgOAOmEMZcZMCLOyQp8I34GbUQqHug02oErM2ZWAer9lLZF2H7k8Q6W9NBz
l+AHfeagBZhwWZZZPitMo5/1Fk5uF0hPOLd2VR4zjvqsVR+IS4WctNgFEey6xAu1
nL9f7jnsFm3tKcneHqgSBxv8/KY49ynEv9rrxbUNKEwbmx2SDzrPenwwtz8gKtTE
5TxSfrvbwp8K2rpFh8adK5KSdhVyazr/ozHpfaUtHDUX4YQZ6WdAg3/UEjOVnUVY
8PCNmgoDISoKFxpcp/W2jmt+gEUF7omK0m/2wURBN/b2wD6XkZr7ah1OQslZXOZ4
w5pm9EJPr4uLXzYIfhzVfgsGrTIEKQBQW1lvM3k59ZftJ+U2lXgIm/L/B4QMvAwb
03FOPzmpf2tJBlEUikuLoY6WyJxlD5QL4EmUCqZuUghgQZg1rHmhwOdjm8htH/Ia
/ykG0U0hnVJvcgDRb0aifb3DOhjAAwacjsyNRq9/rdhRRkLUIOSGivHv4ZO0ICvi
Ze5rgsO3iSnzxi3WOpdoih2L1yf9U0pG2Dxpjqnmu0AJ6/BXahLL6lWB4w8744Ky
bgbXRI6Kx4MCjKJz+Ckz2CPuM1ynMbCb1Gc/C1VkAvDVLISBbzhReY8NSKknCeMB
20yZth5/2ca/Vn0NTm5jkIzq+JGxSJ9ruwhD+RftF3AF6NcojBJ9Mn5SSoR4pp4v
lJAplki9H775nlD91/6d+aRKIEC+j6xMT8x22Bgswn8nKZsbNCzfJ1OBonpHBsK2
XvU8yQFoFGHBi/7FSuf0f1UZbXdOCprUke52IPaSjhRsL6GUPyQ3TRDkGLVZI4xW
rT1RAZKf65whOStNxqs8oKO2bqVAl8ih9MilGT7Id0lwV01vf47cyWYrGcCeUlE9
N28kmCFp75ZM5xZProSDngt9gdavdQjGCvbebg5whFMR/nd0ARkToQDtvsQPKHMa
FUmPTF4O8wpM7yzAIaD6iZy7IZX2csVobBmbFZkM8wmJkHwt+RTekpFah13F8y7F
`protect END_PROTECTED
