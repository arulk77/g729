`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSHs9HYWGQa6TMGvsMJfmQmU/IWuQj5bWlI4Q4X6/1THA
tEA6CS1mfBD1BYu9ksNRe188WxZFt7K3kwZ1DisMyqSza2oUwUoX/SOV5X36hgMo
GuPYCva5M2z75P+M6eXSy1NFobCGDNDeylEHLj0MkQbHnPLWy4ZOgb97frolXpuv
Sxzv7O5ZrPqkK8fCl6+GBEossi9C7GqogZajDdfvlMDDrJZjnis58uTA04Z2s6Lt
pasvs9ircz/e24y7bGPR6Od8Qh0Xi+AOZg4eUAv9eHpQUsDeFEeQu00oL1wa2CFP
`protect END_PROTECTED
