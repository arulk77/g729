`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
y9UPMXUZd6BQrPHMW/O4gG1jrKch8rvIrm8np4Mse+RWYWttd463AkGkecVGOL7/
TtRyb3UZ2xFwuIQUxKpaBrQ4fZYW0puF1SQ+uI/nuXj8qJZG1RR0JFo/ec+ytu7I
UjG8xqkvzw8JfTTQmDqivdqMMrpcsHi6i3M3vK/0FgzC76E8jN+PmbZUIsP8awK/
`protect END_PROTECTED
