`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4y0b1xcCFWYRj54qZ2tsLW5Qql3trPJqVkFfmVwdsgRA
BQCKBYMg9wzABLYLVEktxYayN7Z5Do6bGgzncl7yoVMEM9sq0EIXq7FFbft9nJlz
kafSL6rwoTeZfspYQb/qsD0HhAp2YCRgfGmJQrJ0qVE5bRN7xOTvGCp6Z5x+hJMd
F3Ky1zd6w/rVudYKm6F5wFaKoCF1Kt9N1POuFFfFE7C+LD3EFP/4q53NYDYNNAG7
/H8aUTwtK5j4snMQ+grl5Ks1pxRZ7zi7vWALgj4nWlih4shxCfD1lD97bWyI+Mrp
tQT9MbNY4wB9kwzKschZb8pI3qYlXD4PV5GSksrgJZuCFmrOwGQnWZr1GOhPwhZh
MCIBQkrY6k/JdDJNXwM++EaWvm+ZlX5JWgJnJf9I3MBwEP1ybwLTzTTdR8CFUl8r
e5DM1wcGbNfTFe7g2Gi6wmW7UkdRsKs40WZcbbUMX+4pr0IGY+xqaPTUjn9madeX
ICE1RGwxRIaydV9pDfSMAfPSNCNMaUeHIh5bxZCvjqtrSRxSqFH31wbHogyNGBby
5Rp7RNsUs59p8RzMFQQqIXeBZVjJIfi0ANE+R3+m2yjP4UraKfIOgvG0DZ2OO+M0
f+fwV/eAss6bQa92Neb0swjPdX7zE6pEGNUZ6UMHSu8eGBdZgKN4H6AmhVOBfT7N
nhgiCTlpenRGNb8aWoLa4PDhKZpqVzUjtyP7jluQSC07hkpu4fvFqr3qgP6ZFm25
dWb1plirNbYzuVuyVBxwLq4rtUgIUtpQNbp+rmBjkRJpEb6GO7WXxsNN8UNAoz0V
7aQY/bV/bny3Zn0qdMjVT06ehikKXhNxSho76isWSk6xh9jA0/w7JxLvQPdNMxss
lPmGUSrflISRX2UfGxdh2QRrPyr4fhR1650CNPbKDdEGUmD08hLkNRjbCFcwpglD
/gXYd6wDEfjDJcrRiRMKxtPV5GCtf2O0STmO04lZy6uvJ60ylc44RaRtne6GIOPK
5U1pn5z+gJYmRENSWGRxj6YtsLKNqkWW00d+2L0G9pPZWWB2xntIol5xf5wtFMhs
CUH7qPK9ltAZNxrrTuzqXZFPmUDcTuvbzsneideVFugRp1UFFiAgFplRTQB/fMT3
GuMTDLmsGcv9E9K+aWX6wuabi2haqMGUtHs4P9rsm3uXH7D4zHE0kE/mTmQc83oZ
oQo009umAyNlBDkjoKWaWUp6vJodPSNuB0+ZrXZksAJWyZctCAegLgTbaNY0wCCU
pCS1wYC0dxngr8hZcFcFkdUpCkjpj9YuDAHToqTwyBRaygV2effq6smssUGQsUTy
hmoN6CHxhnw9LbXlk1rJ2OZhSMYyCH8uxQzMkgymzQWc2FTAszDBItVsFW/Z+WZs
SdM9077zNImOg+8m73ABD+o0rX8SRbL08dWTPsq0uNSDbKTV4QNGV3d4R38SVSuk
g4AUIVINOmlilWw+VzCZroVKzEm4J7LN5w6dLz3tzYVSBSu2RNSUtXkJI7SVR369
OVT3xVUeCrhAiEg1vJimcnDeciDZUI6kMy9kU7hS4Zd22o//J+9wYUgufnMTFfZ8
efUHCJEWXd/qO+5FWhtNpqu7+OFQ/QPaoYa2p8qdf8nEuDnr8wTyaxsDOQfKcqSW
bv5LVv7oswyGqpaXvoooUHelv0Mh3THZaew7RC8AAkdlU8MjA3K5j3GLmnnHpQXs
PMCqwTUo3L31XBoQFWUoj9cI10mgEsj5/QwW5zcvqbvrFxcnzNPykoW5NtuRySKI
jDh+93y5ECPAcu0V+ZV4e/lJIA5SkHj3UYlLEQ4k5nZH2Z6m+tmMEoOsf8sBM5Dz
`protect END_PROTECTED
