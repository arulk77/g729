`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEJ71TR/ovMl4w50lia9m5Ejfn2dwX6lEE0Zwfr6Kc5Z
coQngBJhCxwY4pUeO/NukbjjC5Valw1d6QtKc/EKrGsQ/Fioe2GbKRlmVjbq06JC
ucf3A73sMWmCvRnaHFhoPPGknSVEGJA0NyyXwZTS9pGdlTvOaxlugJ/8kfTU3Sw1
ZrcXscfKc9Cs4fAtiWAG4ny3uB4V0CZEBc5SCrsdj/zAGsqwHgJNwr6uKKwt5kg+
t2fR4+kKK7oZ3CDFUDJUdg==
`protect END_PROTECTED
