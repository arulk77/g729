`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/ruOEAbJAcdQKSbLUpchNsJ2w9yDgw0+670oylTD8+K
ppYXV1WNtT0pV74gchgZI+pX+eht74pyNyRMQKv/qefavxuLsCjS+eob02zr0dwh
aTloox8RlkbO0PS6DbX+emUbDo65fqau5W1HD0sRlLx3Mrm4GoSV0kvV/hmARi0u
3trk6Z3yNRcVOt8Hk1oCZzVTjsxMhM2K7S8WzFG6IxLKnJevAYlpTSje08rFTSfV
akIySYiAkyVDi9WLxOuwqlltlbIAgKLm5DBIM4TrKa0=
`protect END_PROTECTED
