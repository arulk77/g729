`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SSVHEVwomBoHEO7leDw323AXrwrBryd9N04KvWeCOmWM
EdFCmXEGUooUb0V+rPM88jv59O+/yavboFg6WW730uhdIldz80WyYZq/wBy7fQoA
v34ERpc+vNpR9SRUnUB+S5DcDfOJo8G5sT/GIr8KYYtecUS++5piib1NgR1s/eqw
yUYIbd27w0NS3j6iAexL8FUTGzZ64WESjueVh5iRpHGd87+TwNhgb+PegRytDD7K
h61RsdWLZOjf0RWjkiZDk0LeFJmtqrcrRDBzu3qog/LWe8rRhrWRYKt1rXzaZxL4
PKx3V/A/mxOLmuDbhCVZCAu/wRjJE0EWoB7JvQSso/TEiZFJ2TRFrHH3x+qTUPCq
zkP9nFP6Jyz2cJfmi4P+j3kRvAxVCaqts+t6wQ7qmoGqUQghAN2e7ysDDcVd90ZL
tZhi3Z5ftN6CdEPilB8Q4QYombxDnPcENJHQb1zdx7kN/8qbN/vyiZToN43n7Q1e
WhikTejwlx6et74NDfvHm3BSoTqTFlifRGcDsK60u/5kRw9oCYPxfCRZIpQmEE8M
n3P1nNvPJU/vT1QF+mVZBruRG1mLA5gPWpneZJ1kDQB6ECpJOJ5obQueXobtm0Im
sGxSeBOaw2B+T+bXyhTqXTqKwZiFQjqCs96iTlEmtaKv/ZypFHblMQKmWaqy+0VP
X8EXxDBDB6vxHVC6B+MKb3hLYV0/0Dwi1nnz1zuo5c6/QppqCXDFtwaBZ9PShsVC
lZnBGocCrBXMifPXCCczFGJvDycZhBva5KdwAma562bQbJP5dbNDSb2hLYPRy6kW
T4ih0DhiH8H/V1uGg+sG7BfKiaYNDVGDI4RUBxiWvLijUOQ1ogAT4DFuS/spDPA2
brLQab4PWcKJsJVYK7fVYPcL1y/4jPlsdD1n1/dE4UhpMeXeAP/IOcBN4wBNqsq3
YIpXAW05/oyLNb/xjRdIyT9519ZrSjwbrEgkYHZ5uQ9gdrAIfUXaGmJrZEjluez7
OTRcufqaqa3G9hNeNn8IlHA4vnfJqHyqFKshKwx0PIJbRlvbP+Th+MpvBhMj5Vvm
f9jB+EpNqF9CFWHq7Q+zdraBfQ41vYTdqW7O0MgQ+q5HnFTAyjVFAvyBE/y6wBuM
jREY7d5e+YZrkGU/K68f5zS9ygKbiTh1Lhkz7eVjxr/ol5Ft7VI8njLaEEDYXPwZ
12blUTLNAjIKh+1tGRbGOg==
`protect END_PROTECTED
