`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TtMjGbuFFuMEIIjG2qjqhABfneJoUr2EpN1LSq8GutJ9xKIKZIAGULbCbzTfnarA
NsJ3oQisnIdogD3uh0RV2p2sXXD0efbe7DGJAnrbSomwaurCFlJYKJph4/74+o7x
eayNCycmxsLI3wBXSmOvbLpfveBID5ON+zCSD3wX+zkQsWnRpT1vXgO3H1hW1/Jj
fr/57CDD9xiRLwfdwZHh9kHxy8CUjVeGsorRe+YgaRJuV9zbIgWDC4FixDR/kRgh
FwSx9YjKERbBpoiYwfCY9Imb+8V3YmKnkMa7n3VCgLwgA1cwJscOFYtUHBu9g5B3
mY/jciNJCgyBuwIeg8GTipQwv8Xjihdfw8b1+sYDEYsl4CEXHA0tjT8NA2BrHcv8
/yeUOiGJUDlzhU1tviMKscyfrRmL7HgMILKv1Oatj5GyqlmmNSf1Z63GSRp6jLro
RQiIQlNycbE4JSQ0jtTzYw==
`protect END_PROTECTED
