`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDsDPgwTSs/R9Uc1QPSgVpG9eMjugDLvYC2pr5R7g8cg
O8h0QnCxDPVGEOWBq+cHl0olUpRUe7+JQwuDymK36evY7bVlnvA1Jw8iIt4dkQan
CBzZ5AoiVJtkEUV10nkYgnZwUeKPzKi5wlH9fmbb+6DlxIPRgpd+tR/476a5BiQc
GHPH7HQQQ7cL3XGfKgvIUUMhjKyAEmj+kDuK0Fyxkw1//9RSMlF91kRrd3CNXBiB
I4lblnCMgohOtfMHSZSSMfDIGTan3Deo6bE+zXK9jVTTU8tBsG5KN9mdXsizXqdA
kxFV/TbBPGB8G3kpmNu0RmNnQgFdrjzF1r5xArRIq4IxC7nG2TceZspScjYMYF0f
7kU7wBu+5tlZPq0nGFjt0CgHTxcqXsZmWIR3tH4Lv0fTf9y4SfGitOENhpZpNi1q
OOc2L4783MEa4D1gFUNe3I4mVFx3DvlJiUtAwsykSuSWhc5hvrg1j4n2mEGmyptz
9J8HaFdva/nBiP6MS7NsrhixNY/L/0aM7VCz8Ko9+fS4Uv3hASQRdt7dSfbZh6Xe
LIAG1XGn290VgN3uNAJTCFLzUlAIap1MmdL4V48QN5zMeM7HIgyfw6rKF91RG0+Y
7vahSxl5sjgvSXMURElMfiEfFLElUH6uN90l75rt0XugPx1WaWhC5MKfDjBNtXq4
78VP6FQZOqdl94kY/foVVYfHAubvfglk97cizNk2PuPYXUiOlY3kDiMmOy0RzCCl
BQpgKcRqKOV3UkUH0sqcxib4MlelXwUbJtXay1+pIBwwLbgknxY4OuiRp/mygri+
z1Cnc5TO7MdjMnt76I0Zj6Q4pGSXfUg+9OSEL/wedjdHHnaNdMuf4FOzMjT/8BOt
SXJdMeARX065dZR20AFO1PrMBV3xrMKENXFBxKOp8WSFa1D4GZcHb8TLGQHq86jI
bhwKEu/R8XWqgJwLkG2HcKygrVE2HmGD56S63344weGgssSML5s16rkgcst+8Ixt
OhnuMxqyxmqXBNHpZCbLFfHZ4/L7TiJmOcA18f1J3tYYunErrkESGTGM03OP439o
hzNJ3EhbGEFqYsHCCSp8OSI4QU87EHgckIRLWCfLandajunxeT43bje94MLfRyyv
hk6JWWmr/ViNWwcJH+rhIyBOD39fPP4F/mF3ovIWHMhaQE4BgIE97CcQpMwka1zF
xAqt1p+NguwpMkTaNoQiAQUH/Nan8va9k4b7pKshxBRQiyDCqCDQup8G2O17U8rL
CKBpECPmJ7viCLHO7V1+nptdhpkYn5wG9ktGHY7Lsatk9AsvExs3XnRmnp4THPul
YRCdgtg5l8VqhZLiECii4fw7wUyCEb6an8QP2Q8hY65JFyRT03A13mWLR06lAx0H
awZvNTYC8/Y5lO/PLYnZmRykf+zHxsn72APwNwT4/5CO/+tmb6PXtc2eQunF5+38
X9B/mMZvAIRZX1yOqECpQTxooNhpNu8h8PEJW1+ZWtGw43YYhAZBiZpL+Xn+wGmh
VujeD1JZL4EPXwVMbUv2odTlcJ62K3gO65lpbYyeSe9doCQO4IqHR3PrO5Fiw85r
TTZzMFDWpGbavoo4+O/OOV7mPCLgtf0bMeq4a8vWgKc7MMx/SXc3wp1jOaEaeZWQ
9TbYk9IsMANB5p8V+28dvwF1slHRzjQ/Sc6JUKCzLyz8BX+SIQ5UFo07Vns39wSK
WGCKKgWSlu4IZJMTDT4zcRXmmWh7S6BY+CGWthVhly+t7Id7LtOp8J5CHHbPn437
qSdyRqkMB/gpwpsPYkXPjLKICP7wNV6DWo39vBI+QiwTV1LfE+cRRl6lA9B9jOfj
c1f/pVQifmglPYy7qY0zxctJWxkpUalhYyyzXOUR4RRGOV2fS4k+zQW3ighJBrlJ
OLyLdIAhMwJUWKiKArpUW2S9qe7qJmIJR/E+V4hk49h46aPrFRonX/ZQecywl7b/
S1XBWa+wRvBlqzDm9lDkBNKIAOdhk4NZ0JeS13mKO7M55a1dkCE5Nq6LWMrWZjYa
B9TFFxCYZ916vxdCUEXBswxk1kbpxtvTlpZSA6vlrvOKARVD3WCFHD9JtQGB0FEN
9P4R/QgWnN2E//nDCnmGAt2YT3AzsHbeCEsPe9NZi60f5FjmqlEq8Y6tDoK/QfHZ
D48eIlQNwzGaTthLeBv8IQ8xISXynS+K8+yj/Yl5MkspKUh46brm9T87/30khM85
z7pCce2PfoOuHbG8r44gZSZhh76DrsNebaJJbPnvZqz0MWPuLq1NxGsOmF9Si4sO
jvt+4flJeKyoaaQKJDlYKQ3cPa19RntidUDqW/C8XJJC44DSMXm6RCgxZ21p1CsO
LZorsO+8cCoThFxDbxyQ7UM5xqTQM943BqPaImeuCvhChoOkUiUle5K/Y50DDs/D
cFOPCbiR8WEaQQPz2ILXiGNA+a3XouQz4I2HZjC+RdP6OWs+23mb2ifHA52329Co
9V1llY3GFr4tO7QuqOfLRT3yQ0bbI8s/vZ8tSoj7Kj5Efd+OhRu1/VDiqBnTAYC1
XxAqHr/LGvIil6d+4inm8iGK+TN3wXHFic7/+HZWF41eqr/VqlHKLt2EUHcTEpW9
30NDsN5jBeHmPhTBiJvNqg++wziUjLS1/SUFlXoafPXIaf0OXVC5qYGMuaaCEO3N
Nqci8E02S2e98E9Cyd3Y4LH8P5B52F4enQMNPcltax+W3Vk6OxvbuUDRRz+4mtUH
kqljafUYW/rCB9aiTvTqh/TbXtkkRGnLSDCMSjj0NiCZpXHWYgwrXCrJB7wMiOU1
oHjuh4zeIlxhNe/JULCcr3988DKk2q41uGAnA+5x1F1uH2gw1+sx2HXmuMw+grs1
u6XVftmRPU60XQINLdXixGYhJmRTP5bASYLJUNJBETQsfaaZTsaR7BxHBUxM7BdL
rZOr+6CyQdw19tDheAE8oinOgq7za992Sk5M52ym4fL/lycWsZET0iXNi6rjLoSc
LK3T6pxFH2wq2a6wFj4CEYgbzsn4ULqz7UjeGehFL/sMZRFDXDSXxNk4rNv0QTH8
vKWOIJ2aptg19lt3QGHpFv29+b6mfBO3IJnBH4gxqM5e9OzSMRphuWqJjJHmDlZ+
jgJb674g43KcTDxHwu6HKXwbgqVGi73y1LRyzpjpftOESDGJs0eix6BlbnWP7MJ2
GLCBTAbe/zxKqJtqMuRZUFa1yv4pqJ2WgJXsGDYeUPNSnqQGWG2teInrsUUloswf
91p82MHn14cXdFultKzMTSefmQIWIO/5D/QHqR8pgMxopwakYejXIJ5oH9nAcQTu
L/VtLuwRj81GjNYIoiSO2if2ukbyxu57X0Ws0SVKGIFF9fxALgB+CgImGJW7Votd
uodhxtFb/yMGINDKr0XEcNp/QnAUAb38owLh6few68UlUBqkOv7iEpb7TH64bV+U
oFyRI0LlJ1XOy+ZVENzoEtuq8nMMzd6l6/44lKuwyBU5K6wUQ+KYFic/fSGx4txr
3uNaiMYmV/mdABo0VSrLylD7EvRymTXoELLQB4bbmsq+EUgFZl1rE9l8bpAB6QJx
ftmM7KWtnRCghStXbyW86MIDwCo8lDq0K+jvWo85J9GUq94t2tTZh9nXtKRbfJKy
MaCF5YyLLWs7ji87t989ZkZfX6v2/fIaBWI/jQlRDfJbIobj0FPKg83kwcwhrZe6
1vzUCgnlxAoi2aVl6fdYaHqhUG1UNbGKsubex7ZEioesimnmjOsBL9XI2q1ZrOUa
4/TnLM7HUZ6u67nBHWhAyz2e0NL9pNtmMDlCb4d7VcrDE+8YrYzTWvbdTvQ6Tw/p
ysHkLE8HyaF6Fe0s29raErkNF3lz8eqvR3BsIi4lg9qSQ5cwrP+LHHZPVx9upqd8
qQJfGrm/1eTViwKZblf/uoUdtbF6vuzx6Jl3rnJYCM/Fe4NrH7hXngE4ymTM2TC/
5QTp6NfI28qDo+ziWUDunFo79tkoxQdy5KcjXhVvcPGuX6q0hS1+1cOc/3xZRnuQ
Q65Oh7dVLCaMESwoRFCQHKuhSpQDLXZ59eWXuZBkA0juFtS4/lQNQB2c5nXIrwVK
TmF0paHIO7GNwuMmCvvjferYw+qH66K7WcUJyqb7uW1TjyQq3ZGtCKuCcLEajiqn
/aMJwxPuNb5kR6W96wb+XF2wLmy5R2uMqaPzZsgA2zXIX30JVUwK7JfaN3afz9S+
XvfRzxIEBGQ5GMi09BMGgR4HJGlyIung59pB8Q+ilWMGwv12fDs35a1HnyV986Iz
lPSA9uwm7Xd7lRdm9k7/rgzVXXyVCrokr7J8p4shPxRzXOxrKvEoD5Indd4+zFSR
epjM9MZ1Ssr+VD0BemS6jH+S786RQQmlFND4XXA8HgQJPM+aQPKmdck0f6X0IvK0
ZjyDIntNr5uiEBPdtx0mzT8LQ8xQSM26SaBrQhXCoWGIhgqHbnXDXgnQJZ9XwErq
VOmDG18gsCdrtIW2urP4Og8Pjr20eCLAj8g1lxi6Ro4P5rs6Y6kXaXdUPMlcvN+q
DWu1VAfmpRxr/yUE0CKcDzhQQmbHZyivo0UDNs9gFRwOM/aa1g24qCI3P19+tkBf
0fU+N3S8RMO7cflGmSPPKxY77PVjXYXAKvOmLUXWFxc+PaZ4JKJDKve6+xb3hiG5
EE9uorkdvQy7lxWH1ss9crTh1P3S6iUapGri2zG/8VGSbpHMXLHXJdJ6LZqBd4o/
JP79azZTlFnA7n7s1q8SMRqBtvQFnAOBfyc7w728qgiIoVQ2B8+LzXnDPNR2nfXX
r4tkCfmUceY3+zKXTE/AJ+opeX/E3x0LWNOtcve75bOTF2cUdFydIW/pEBrPQPsQ
2+P93q3c8Vdho9rvkDKAybeCMYeNeyvcAyCtmYVk2LpLkMHAlrbUFiEL/r67WX6n
k+sWpIc0w0/+/cguPthiEQJaxE123nneAWsWF2jQsuAEjcE5MvDebF37+d3yH9Wn
1NXW/wvPD1jJyKcvG6c2c0dE7AR7JDFXu3fftFVE21otpkLSn6E2kzeOhFdiSdB8
XBx9iaPX+gh1GNkR+oLhEfNotZFfXw8BKLHNpmKWsQUt+yH1DyNIoYTYm7svHwtr
3T4E4o8cqjdedK/liMfKplX9memkgKSD+CzLksi/yovpbmLrMFeCU0jNiS7tZ3in
dS7aOplp9d301tJiAsMqcu5jA8MTZjcQf09MhKRrMkqWVeYhTUwrwRq6nVCDK2lt
k9GecgyTaEX/ipEUXhM/na12ULzvpBXo6xdjXWDbXBinB0w1ZyAJMncFwU20bp5M
2z2PPmoN6T9BaYVQoQgfHfeDO2vy1IBXcU5r+LUsHgZGYVdGQBUpzXDz2US5RuQN
yIf0/ImmaIDyrQpnaoT5+0/pluffGysqtDJUfYeOOC9G3pGmKy20jes/zdUWlzJ7
kHiF6iHDywFyhllRSIdRFe5MwOFHp42hhwRNA+XUG7wpAcEtcmM9OeMCerAb7kp9
4/m5TXpnr44EA4lKZnajyIFYzWqdXlThz1CWMM92JnG0IxEc80QLrY/ROdcaYMTx
mc1P0/VrvdU4c2fRwyQpuWxQsI+1f4Rt9kQqeqRHFHF0AxKiidrJaGnyTaW8n6Vw
sPCrNr8PIH1QYDuOSjVcEvkyYqhhyW0XZmEvHQkCMZR8U5t8ndJkXZtOo0qRX2cL
03h/CU+F1bjVE93YpiehP6uMt7EWUNB/ns3i84PWWkj1ESZRbr9iOWOGxZ6WYPeg
tZPueNk7lMAecRcroRPKcpg4MDg+M+ZTA4czuQAYQlTy22AxU2Bjn7K8D1DX0uab
tuW0gLGF1Byo7TxmuYxanu0S4xIWV2MmNy3nW3MbMPQQ1WwN2uCrI2eH+vDLqqY7
OSHIkEjq5FswWlWpLPAyMAQVC0p/bSE8zqjCpykURiedDWTGgZ0NIjSrEE2L5C/w
IcICYR5IsH6wNTLkMVNCP7zJb8XrosRZ9wkm+iAxa2isXtGxibeYaO4B/qIBIuY2
oLt0S2Nqplnu4RSRQehkKwtpZiSkNUfrDYlOw5mintgQTsBNGT0mvs/p0uuSbMfB
Jrryn3GGBZCS0UAj2q5Sl9Pm9zGgYwUcS8h+pMyK1kwU7wuE6wucTW+NgoGuVa11
vzq2pzI1hYLnea5cV54AiYg1gNyPTRxKlUw2TLq+8oEuEay9BrhCpM3e7t92RbL1
1kRjEWl0yfpp8oQqEvjxC0OeXH/bYGhllCA19duytgQw8aoQ/EWf9ImLCLa4wU01
aRNKdFTnCSlINfgFPhxhQrSEtbZFLCEmegzhM00wkakXGjBfZeTt8UQJskWPKoTE
Xo471B//wKI5odJEGDfhp4ROkzBCPsxA5ppWCCmxU5+g71rzk7Prpuo3ZIjmXZxJ
FtY1ZIjoOpK314JroYgQ/7qbyGUStrP2K0bWjzLRCV1F/Pt6J05f78xLR7cfZVur
2bJWyzHmaIb1i0uR30YJcV5ghjQdQwo6Fn5dW6j/azJu6l36rfp0XaC2ZhwIRhEM
lEoTmStn17H+lGeygAmNPPuMbRZm9pzlKsIXExBFPvmMi/gh1kGg/7kHOhwbxRBI
P0iVGQhmFIMESnf0HIQHGPXDxi0vat5zNZaZ+229pLk6wqhyD+6Jj1anY5F4oOzC
bOOTezCBAj5abpXZXF+yJCGadLGt9qVm/afaztCoVQmBVyPjUaaOr1MvWtC2Pomf
iTKUTv8lb4zBYXcHq0x76ztmKiwKT6AZHCp3gOnvuSr9RlaPsDaW89nb+iaP0V+G
DHb7T2zX7HEj4JAUmbh19OUmb5bJyistvAZnIHtTHb+8HMbER+sw1apgwAjippUb
yPgu/GddSuGWSIIEYljKYMJA/PZpQ6Ssxd+8ODoh9Sufp2D/bkTbRfFE69+OYgA3
YGroB2k9zOYWlFhpm7JfYSc0lrG2pxlWgAgSsKVHDrw/4+fLfmanPSolxHhGBEdr
rXHRyDx0is/9F8U9ph+fV6U42Vhk2qEschSuj6dSJoy/MvlZ2ICsyWB7a3wNPmiD
ogc2K2MzSBDIe93wHpowo8p8XxjMdmsvEM5bR517kysAS+se7WdVgkFZBINfKj/c
sTNz5VgOK4J+RGT8au4Ytm1xhFN9FMe0W45MBPo9gsLbufep/pS41hHETce3GVMb
5FC/4d6ztbhLGYPbndkBBWNpD9/P73bJvHWc6cPSUMJkvavS48M50hCRsJKde94D
0O5lftFF+xl4mhSCl8tkSJQo9XJ2upB5BqBBbpN2BoQhbYOayMTnJfYp6w21ohWg
m1T/gWWISdlLAsP9GwnnfpcW0tV5tCmUjZm+PEe0PpWhJtKGW4HYGFNtIM6vlYOi
puJA3Hz18RMW/BhoOwJcdiP0NxdDy7VH3zl+TAtR4osgXl3elU4tdLhmqIuuzimq
TB18US62olzLTr4l1RIPWDsDoxncmBfUOx67aOq1xUfIglM39RK5Pb4ZPPt68QMD
dkrsTbfKfI7yj9Rvhlg+6vog6ZKLbvmyDPNuvxnX1/bWFeoLpv07VXns5lLCWM06
8nqi7fBVxC1wzfMBjjGE/JpbA2XbuCcvc4zz3vYA/a19LT7QYAwS/sr8fsjZyeBO
mvLLtkUICYpIShuBTqUvIrSseUnkDGKt+DKM5DEE/0RPt0fDOMwdg/ovmSzr8C9n
4fCmW/hU38kdW4ITJZSkPfDyn+TnPEqT4+mxx06ek/ejRppTrqW0Sgk12cz9B9CU
0CjWQRn8pztu8mWCc2I+9NFF2GMAGaY1FhdsfKXVDXxRkixVHfvZnv3v48469Mx6
Bl0KsDuo6KQdPmgfMijJ4hWEBfOzsKgHchnNXuBqVFeeNMlQpRZz8TowKSQmEkrO
/t47hS+Ej5OBeRFPWE6jJgm4sKAexLo9aPOEsCVMH7Vj/poIBVJI90eTY5IdOcQc
5d75CTdbWary5PC+jt44e3eK0zcdO2K/F22bi8Pr5doqcgnMy7VqNCFjtOpSmzA3
9YKyLBIe1hLs2xbsot5XDJVSJ6oUW9llF+wnlBn4yFXlslgsqVl1Lydk5pKOzEu3
q1c1NNgmIiyrBXAduoFizgQmEcOKkH4fYsPT/RKeXmU4BZdqOoz7YfZzms4yDAb1
Cejfri583XTuEIYvoeCB23jjJfFEgUI7vK1Jfc8nMHZlBKEDjhp/ebxtTkKG2b0T
56TknCsCHDOFhNoEbq+CeEjRmNyMXYBUgC7R6F7pVJdDGWXUtimqEtOt1AuI2OGS
aHsv8a2KAK7k1m6j6u4Qg4BxFjK85A7J6w8ClUlsmmrCq9rrtBh8E+LtkIDpEUK9
fzj0/QjeHqEDjtPtRc74Oo4k5/FSvuHhYAe/7i44dsZpaSu/9/nx5DyNDnIk/t5r
1KoTXNUcoHHBoWH4Sgw1z81+JKbkR3GVzqRSIraMd3aajKteLSRPDFjJjy30vItJ
qFmwaPQwrZgV1K8JmxVVM+aKKYqEc7yg8CfEteoi/RtvctM0NJ1vykv7D/Iflgbp
QiAfPG/TBLgyUZ6uM29DPJi9N8cZffNqoC1EPiu+EXIv8K7m9hPL+T1kI6vK3d+e
CQ9wplaKCNMS3zKTLL/Sq6Ci4rjCq9OBzT+x8PINN3d6jjrFxXyhH+UVdzzjmrc8
C07+R+4nXbNSqhMztSmSX6eKd4etAf3du8niA38jjuv6GbItpcekepOIQj2jRFrW
qgklwIBbOIAIv82P4Qv3s3gWoqcdRF1JGM6EQ0xlRUflyoBa81+uMvwreIzIPUvS
Hixt0/ncxJAq9PQL0nKLMZtMGJhR2mNcJ/54EP5A1RmZwQyE251IkpEK8tqNcYdR
4o6zZi1Ub66sp6sxl5YOFBdvxVriP382rx4Hju/lATRWMJp9X1mIShQU7Af4VhHj
eoeV2S2jZ7Koa9sZPzN4kp+nsLyFSCMnFWr1FVb7nM3c6OEitsqqDteFfnsz790X
t3zNnPGyXHIOhKPjhjNlP4UhfveBPBOE/VTLXH80JJomONXMm2s7vSnWQuAowp5T
7qDcO6yUrueGflSdN36uDvd06jmxC+cfCEUeTVsx2RAnj349snqUpWAckBtAJZjS
wd4mp2uL7BLJhI+0RgPLuq9Tf5/Q1joeu6TZHBEaQiuOWehaFIpsCw8RDfsVnwGl
GVXhn6leBKNcu1u2VaQHUA++v8tnd6lXMkv4tr2YvY6UvpajcoGBeH4x1JBUnHFS
NBoHyr/7CIINDKd6Qbb6UQ4Zk5k/iU5iKdJw45171lKIZ2jJ/oT/uzF4lUUuDyHc
uV5RCi64GKE0heBXE6KEaj2/YRAtyBnXANeYCMzjlW1fHIJQBXdwH6WrnUTGcOUa
OijpmDaxVJ5I+NtuyzhesL1uq8qIquXOu2cIiTTv8hXO5UaZN0ItVSF+altwqA++
9x+cB3ueCBIVCQ7TZ55UXlLk9cShPCqX1ZjLHMDEtF4r+nmknhevw2vgo65Tv02w
Fwd7rHsTdiDUB2edDgCU6p5QJq6G21wGJd4hUqwC1HKLqzlzMHZA8VGruIVV85eC
g3qKQGtS9aB/osRGUstpqk6PLHUiLRtjwkiiiosJmMXHfzxyIYh6m1zK7fIXRziV
OihqdQYok7cShyS4/330USoPqoV3H8Cg8sydcDx5xIaapHwhW4hthoHkxZ2jJ1ZA
EjDP5LWD3oVDgoVEYKmeo4leSYDsL3j32tfUXCeTojJKJdogaB6xTORQ/Cz3Rh4m
UeOLOSwUXu19xO+QuyrxGs5f5s1tPu3aUtvr7hjMi5VD2qMtPr2mG0Jd49f0lRXc
eXTplkNqigVIF/6TIwdVo94WPs9nJ7mS2DTBKJWOYkXI/qW38pYzbBWum3iGX4/y
AedAUpy1LnB60UpYHhMX0JP+TE9yMHFCDFiMHuasxf5JnWdS2VDmCk6JKdW4+U1s
U5Sfz5dZe5qMtKxnIE3RT15ovk1D0AQYc2INnjgBiErhDdEFs83GvgXx+mGIromt
4rSFzn4H6v7nkWnFe+aYacYr53LUCegXdCqQHd9yXE3qCRefW3tdxokYLgC3nJDd
/u1FlRU/awVuRIhhhbAdrn+zIS5hnbnB8IxuTf8gEaU4fZLZgr8MjSXsSygHzD7b
Sg8jhDktQ6mcHYG3Os4uJ6gUT+aZKNasRxv2mJIU0n5KWTvwKBJM3szYM9CcgJQT
WJGufqRH8BPchiBmgn1bJP3Rn/w80BNNm5utODb/88YEXurN1lH66UX+nY0Oeig9
vtjflNZy61XHrhnu5raN37zTWnQOg5eUWm/QSEuUFDtUb2uFoHGnIGwqaIVFwJ9y
l1+Hf+7tWV3d6yn/saj97uIer7QpT4/yTq3bOb0S99i1wgmrAfKHnSq0RxUcUhnD
MjLKfxW4HoHlgoKkz5NXPG/oUa2BTEYMt/BTR6SqCvzRcarOQQyBTIF9iYM0rbXB
xOl3HhzQmX/iknpPT+UJlsInTYk6C5yvRJDpFNbGvhqFMitXjBHtSl6/KOYBRwY+
gEETk+lSasuo0F9P4ACb6A51YSb9irpHZlazXgcwWP/+B61GEY+T6lG12wZkHyBC
oAMEEf1A3Mbt7Z4tKRpB6bq1lFOHam5zNfBzINH8UVM5VkoEJdIPgeTgid7Kp2w9
edrPMYySYLMIW/O4cDLC6EJByxXyrPGuqc1KbMGG0ruXlp136h0hq6gnDdcv1W8v
/WKyvZRbHefZx/+9nTf7O5vQF1dsjbkcmgEweQtAC7h1FOP3nzwI1YfJydmftgHe
In6GkrBaBmOpClekz08pyMeX0ur104TeDtt7xBEQZ4tASbID0vBNykBKPaO9u2+M
J9NIwCJcUK1JQ/sUzQwfhqNCJKecibMa/5guMkdHekQqj5VLyVzSD9AIUYheNVUk
lCJe+UJNyfrLspbnHBmdX+4W+ng7chaioP6QCUs3YoJzNYig1f7bozqC6doVwWmS
7x0hSIIT/zifZE6JMYwWwx5Jnaxa0uOl39MD1V/SsQP+IvnlCLRadtT7OhqLw3ZK
vH8u1weQF6Z65CLydjuH3M08VGTtOC5fifbsA6VpIaFUqi2nXbRPoTQSM83EkxYr
jSPcApgTSp+FcoRCTpRuHoaVSOEft5AKp4Ymf1e770E0osDo7ncqfBW1YH6Fvymu
JlUUhsQcbDP0CvJUyaPYMkxVLAzhVCJYZxw00s2Edp4AO1IYF5TRDIYBqO/vllb0
NtUIuzIbDUvHwaPCof6HX57No7um8FxB7kQiMhqgyizQLFV8679Mq5CvovcKdi+z
jGi2jraIxfi2H6HoHtpVkT5ZvuPf4HIxV+v5OXIk9dX+sYw6q7CJ9kWm/HdzmyFj
7EWUnCU54bMmqNDk+TrqTbUDbGmMqeF+epXXXXA7tLOWjSDIDk/8jXR8E9FeK2k3
zDExPvR1Q24gKNS6K66dQpE64MEHaRJAWWgn8krO93EedMGYqI48CzGH7yZzij3t
l1edgaR/A9FIg5XvFrLLmaGLDQ38KwtDLyfkkI4gHYtmPBVDvJ+zmK/wLWt2vKYz
cWsdyAs11OAG4pHCIA2kZvxDJELQE7g2MwvkimJSkob9yQHT4cD+rIgDE+l+1fo0
Os06B2++n70UHCKdI9L0S1KYk5vJh5Y/WVGBv/HGQ8MDBgpwECB2avblZjOgQch2
CZGlPdqOC4dl6ccuOrLvSbChzsdVQnQaSBpi4YjvpHS6Cr+Wxid8DhVt4gqdXVVo
kwcjkWcaunz210xT5M3RnCi3bo9ASJblFTnaVN5jJJ/7SnrKP6WOZf6ycEKC2P0S
FNzSB/OxyVnGY5YKItj+ud/z/dGxwykqCZg9C3M6TwwWkk1RIeZ5dzOJOK8i1ugo
wHpV+gPTX+nttlbEO0z3hYuIf8PlWTFs/2xp76472xWfO8mZTGvhckIWW4eeX6Ur
JnJxXd7SWh7kR9dSSf6Wy/YlDuzSn6Sx38pAwGPfSgVJ61NRfuXH1xuDEFDDf1ov
GOpxzTWF3RDOBZavabYDhQQIRFN1qbT/qjXxzE5xL2NnvKPzdVk6DisAOigTODW1
5sAFbaDbZMBRkIhO8AXEhrVsFIaLcO4FXPj0PNgVHr20E51i0GouJAoImvpTJSP5
JE+DITp53lZLTw98jp//201XP58zsrsOvLW+2o9tcrVdXCEFjt95hZ8Z9gOp8PnU
En3pSNSDeLsPJTsxsjXtS0lPHrGMY2YaAeSDHm9oE74S8swq9ZiEkIrxldDM1zyH
GCpAzRSd0HdLXnIGlu3fNdkpOcB7dpnKwJtexuwJipeZjR3r/lmjBNU84ku8glWV
7iKTwEwIlo33OW25t1RvO1g/EE7GuVMRiuhMCd9lli7moPwPR5Dlfi3xZCJPrQKy
2/iou+gR6ekAE9J1QOd+Ycg+DLhKZRNM0j3gNegJpGlaqLC/LfE0FGSQg2LDy4DK
dlb/tN5nVg+/ZOvqW5txf3bYw6AxWVTt5VlHJ6NL+n49uJevNw2dpPmxA5e6kbuR
MEa6vYlEaB3z8/ELi0QUML5M0r3jWeve5X9vrbsJCItbBZwCHlbCJH6tfTBR3Meu
GuIlkGguDnrlMwZ4CjjiUTL2GIK9JpNfgMoQudCFBOan7kzqE7LK4m0PHe6A241r
Q4vNGqjxoYafVu1tVFUATs+FudsDphlodcAJyn3T2CYdX+BjmOKeMNklZFTblWqr
Vfqb19OxqI0/BO2E5BCOD6xU5AYfQqkpCemHsp3aius+6FILxNpuDDbsB3WCxL5r
OIxoH3L7RMSdHXA2ip1vnqJv1IYiibFJ+puYYr7yGtVcVAPFmkofFyi9OC0gZ9LR
ypZzzdbRXPx7S425r3Yk1DQmgtSTLGskD1zjnQONj67zG6/+C0FY8dO19joy8eLs
h/xK9J17DpktX31p4NLt0UNnqiTEkst6pBuqiNzuymwjReps4kRBlRTU83TNyWe2
+/POdG4m7qd+OGU0ZcDPjF0pk8du3vcnsjg1Vu6bBgHSs4M7xWkaIgXYKc8wUwpp
d9CRS5ZwkD8BUWAHFxJdBINIvlQB44JhD+1l4IoA81X6G3GfXMTRA0MOHSyOIgeB
RspAG3GzI2cf74I3UWKFcv1tyTEh1h5AKG67CBb5nJg4YZ4SxIoGFCHm8z76cjLd
8V1nqA4ZVScdyES/U2uZ+LxLrseUEQG++/xIRJHBztSv+jLOkmtXdwANTf3tC9Ns
YT9G2O/3vSmay6iC/lG076Dn3ZVctT98WytoV1rT78/ExONt5iOoIwhAtQo3o/uJ
sgs8qulkrc/J2ixndWeGY8D8aX7jvefxndfz93MMR3g=
`protect END_PROTECTED
