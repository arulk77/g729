`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3ON6twM0bRyFDJLDX3TyepArPU6lhkqWxOspCYPJ/PFq8n+ZsoQzXe24m3qDZqKk
r+t/X7ba7wWhhm2DtDcsKw0qki3X05i31NbSh1LvlhsVCKOiv61F7z1JG0pZgVx0
5aOvwbaustfQsCTWnxbNWvcyjceNZSSG5DfMs99nxXBJpd+3cL/Kz23BEwLG0+t0
1HSDgT1bKlZCzdpxub3dIQ==
`protect END_PROTECTED
