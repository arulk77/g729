`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yCwFUS6gtKXUDDCa5bGH952cuhaFcWLyRyko+0kOm11
9gQXPSUFvwSbw/NU9dETwiXi9GFcEd4v/gYjBBEcA8ivq1rYdIxWYu598th05PK/
MMNZT2luO3j8oJ2Zy6g5yZkdRoxMwv8DisUfu9vLRu93e4Uzz3nQMVkTYwGt1abz
Dlu/6IFk2KE8G6FqiXrbPXZchw/xvx2kEFQS9rBeAd11FNwXl8a/lvHozm/RBZCj
JRVE/1eQXJ2YXbPdAiBDQ+j955KQWG/luypRaKjyMlkjINyjJA2cAIS7Wwc1vSD/
oxSvYjIZtRGIDRBI7nSh/w==
`protect END_PROTECTED
