`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+T53dEcKibSXgDj/8T6OzkGEEsu2IG65z9UB/BefAtj
OLtX5Z4oNvUwDw7RPMy4uw2iaZO+ugZDQbwxDyRNbc5Li7oEPL8Kvq7LX1M+G66v
yU86ulZws2t255t4zeZjMVRQsV4vM5yXiYDXxj6Lxr8sMMBSyPbFpmzzfv4IiD6I
TTSGI23PfOfsz5qqTvOx9R90DADS4HLH/3HIVEp39qbvzlli0kWeUcMPdHGk/LL0
ulXQgHfhCuHJAr5wQnxgKMrnjeb4Cld7Ks50Yvb+ca4IPus68mDLTrLQvPPK1heD
eTVe/CDwc2U75lTx/+PRrJvcIAzekyooT163/MLBNe77hFfnokpQ2/L8E4tS5GSf
/Xqo/kFFDi/yiKLcQ6sLJw==
`protect END_PROTECTED
