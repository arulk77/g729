`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLLB8xh0Ak0zSxFxapcq+DMVAmuUnyTjYlwIl2x6xts8
znkRY4z+hFE+B/pagV8x3/54LzjFfT8Olz/Ux+O5PFZJ3y5pNlCX9vbv2UekcYph
q88XYw6sB3lso4QYm6vqWNRvozN8j1BMvgN8Zh00mJb1EDohi8LnuMOATv/LNaZg
9lQuVVRjEh+l6syq2wbDOAq1cHKt1BP9261c94QHsmw1GtwVWkk68dI34bKoV6u+
Bz/EE8nBK+qArME1TPPSo/zRImgbquF1Bf0rnZZO3SCLmgEbfNpgqTWa8gUwHeTu
+VQG23g5zBLkGJ+HC0k+J8Pu9Fu9+PXDhFlK1OzB6uCZzrfAZELDVxJ51/lK5Nvp
KGJ/jAMHsMH/HrpYUJzY6Q54WVDjkUrTzXHhgWUR+2xq0Fn6yFKrXCxBXV2P4CUn
LzcFPK1Rr376WA5Eb7syml6et5io428TbRfj8+6Q2nnRl24H9RGKnorEvVZAoaO5
qwFXlwHMuJsv30OdwUolrHAQuxSBQMUh0zys4Q75wXmcYs2EktTkwSOONYa48kcn
SY1U6QnkwieTk0RwNFnHhQ==
`protect END_PROTECTED
