`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Bh3Lcpg7q/aomG8aZCJL3+JE8uQ023hnwGvSwn0kKikjh5CvlQR8ljzWxMTUz5X7
U/VTbYCb1wtz81Dz7iDeE0TxlBb/BOAYx9DUVJHnfvg4EmfF1Fs1LvcczOAz7+MB
gx3ueopNl3gDEflfAniYtIsHArcNB7qpsPX0id4NZBq26FMljm/B3eeQa9m2MnFX
57y4FVNBR+J53nf5U6RWKMpFnQ/2Vdek3WFafs4pPAAd6TJ6dW12km5WanDf52w4
NqPbMVEQMWC8HPvAJfTfIkVm2we5W4qUtDG/FiADASUID7tcTvlItOOoBPEU5ghM
4UN+6B8+AbrSi6dXr6v9XQ4hOhb0DhBrAZu2sIDSUWuUKHjT1sSn1sBwOt+KtrHf
sd2jqdvHyN8XrzuTZME6G6YimOG0q+gFQnOkn0Htnjeu5rELFifWWxaKi64o6qis
E8ehjNO0FxC+rnafO2iXhO7RirjEC8xpcElKwO90kBWbyOl4boZKOdtUzARC7kNQ
TSLXHEgqvrJ8I6YRorswk1BjXrWs+mNUBTfcdh8vDlJtC6hbY9mYZXJ1LIkNLQpx
M3GgVrRburY+0IkcVxT+Tf6CPNhZ0E9o9VMTOiM15XvMFx5bJ0sYZKV5sC8+0ZxP
zcK2CUp09XOU0JRpGbLRSb0kvKTQqhrktKiFcbZpN3/H+P4XLnbKTjx7VInmTWTR
tMHh7s8LgcuVxyNRisXBjwIaAsI1VxgQK6KE3qz4QoQxAuo7Ur2Y1Ywh4UvP5/6X
dgv3K2NOKcf2nuDdwNQPb31mUXPizb4s48Zh6vJjTAZGvtLv2dJ7BrVMuaU5+vzU
TO0f5VT+mHqvSHoQiXLkoNU4YmpI8KDC2Y/hhvGfx+rYzKTw3xWgBwL+BGk254Ta
E+MghNvUrnGnfqAlWiogwxhH4kMwuxz7MqN0ATlq5Ck3QFzv+zJJdekKnSXB+TaR
j5QdPl8XZp6ZweoanAiq8c9BHaLaTpMxD+U+wDy7Rc3q/5j9dLwfj0hwLPF5uyaa
9LF/vmq1WHfnURS1vA48QroDaP8NntxuQikB6N6vIlq5WL+OuuDTxCDE3olbCS7j
TxBQkKVc28HzYhpEvjZ05x7hUGjeYlEqzdYvQSf6zMAWIi8rI+3ESHgUgtC73BFn
EgeILLVw4slObaGbhpmX1el7K9yep9GTFwK71Gdy94Dw1XFkBvg/YfJnsqzg+vPn
GAiK6hVYygfbs5lSz+EulfF8VyDUjI1JDVWFtFm+HJOJPgZnIydFeolXDdNbOLx2
7ovSDUWZTwcnvN/q+3+CxguZiKTHiabxcUWNdyw0N2SFEPR+iEkO/9HIG/6nYEFC
jKrFksoDsPVrzzmZIsCrtJb234DDcb3CleGcjHIBTIW5UetJy28+jdH34AFEN9+C
VAcDNYj5C57lXQtYQQM000MXi4aXLQK0AMTYMaxaCeuebIa4GJWYbgo90XLKHdiR
CMl7o7yR57wQKhqKv6z9ehRhUWJTQIjkCUfzfMb1wczcsCXEF+UCnxLtmnpLvCCC
8kvbOQfqewvcquzoivy4YLrVjHjn2/Ao6bxXPCI0F+n4OwBxA4eY32/c03jASZob
r4Zg7oGzgPLE2AJ1D9kwPeXxxwBEaskM7LVaBMek208xKjpfKiJ/I6nU2RoqJcEc
Ax8YRNk0hPgIB1FrMqSU13S3yp6nCMKrTtOauUc8XG5MaNs+RGzs9f+3Ka3KgiGF
EKQbHrvBB+7r1jsclpEXCtjz47MBp9W2ZnGdaclrWF7VRVjx6O05p5hWWw5X8rMS
5PXcZkdSPnwHAzMIC+cfrxAIfQe5FfpGnKOUFmrryTfXLbSepSlisG1YJ6WAujwb
3KI4IQYfEvXQSRS1VrrB842EjqOmw4B8YTckhaZqAOA+H2QAKlpU+YUfnxDNcP2a
EogxZ+G0IH7ImZyIhGewdNnkC2lM7D3Ooe6rWd308PsHPThdQQW/KbLkKtTc4hUW
OV9T/8r4NPS84NN1kU2g2O/QTByLErOZSoQizPldTwLjb7UJndCq1n+o5NIx/s/y
y6G/7HRbqfuRf5iQsHiJhHhybOx4vb7tnRerf/7t2Cy8DHd54oO6s8sxxK0BLi/r
/C0IHfJQ9fok6TUeMrguwfGkEr3DwPH9Ak/FgH4Yko11V4vPfz2Z7JYFscKs8/Z8
da7vTEZsJxy7A3PI5GKSr5z/WL2EiZHGTjOMpM6E+CORrHcRwnhqcbyP0AyxFsS3
kN2NIjV64wcTta8yoVniFN5XpbQsS/KKKi8q6XY/ijveWiQPzFi0MHYJE+hcxT5p
CiqmhrQGPsFo1P0iZM8YFwprGh0bU5M/MWsTgkta09J6yfEYdUK2WVJHcRnr+vMp
`protect END_PROTECTED
