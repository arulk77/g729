`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOQLltGTDCxK8V9znrEoEqgO0LB9Pqlm+RLMykqZ39Bf
Z133XXIRVsOgclW15q+X96V6Ubiy+rpAptWYdygjWUCL2GydVVezX3PvKipc2jYP
ZpV/gtpOq8fqpabfYq12GuYCbWIyC0p8yELVcWsOynmwg2CIda4EE43kUwW5fDAB
XDw42E9pYE8bteGpC2abNLQixfAS5EdCI5Tl31W4nkVcDHnlrnPSvJgj9qn67WvN
wpXrggV90kAt6jFzBsxmdl8WpaLDsUtSp4Mr6JSvlXv5WqS420l/2szE6NWr/TFq
bt9GwwGI89tOjlM4OrAyhA==
`protect END_PROTECTED
