`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
o3C0YDTbWJOdsXPqHE7BrwEwZLf5Z64HfgkSTd49Vl64UGMK7+WsCK2ua3VATCmV
GH9069oxGCcRiZPBas1lr/KW5MwSyxR/N3LxpiwkIyzvYvXBBs+R9M0qhk2Rq7Q/
8bBPyNmdEfPg0nDb0a8gyDsC4aUFVbguxoR9zvBWKpCaltdsmKrN2/DjY4eIdQfX
sDEOBduJtprmwEq6X8h5iAJku8iHyKKVIhDYpw2FFGqdpVLmL/MRmfjuG0krZln9
S0ue0FbXn+nw4+Z3AH18dRp8JsC7G1j3PfFjsEAB6fY=
`protect END_PROTECTED
