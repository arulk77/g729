`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP714IIAua9XFB3HodXEYK6eW0Lyht5UjbfIHzD09YQi
HdETgH28c9N4dgpDn4+HEZJdSZBkZnTD050igXO6dJM0wy2UmWg82Gah3U0IIbfU
Fhqn4Kaf6VpAjdP/YyY9vXwlbIMuBgjptCvVvQLc5pbT/qzqHk1WCWS+obQSFic7
tWfOaiqun8+XoC56prOnVBynRnxAUKdQga/7mNG2WywV0hpGE+v9TdcJSx1fjB3t
TpnMSrCuapIv24LxPVllpDcgZQX4p1rYoZYnXwnaACPrlKyRHFNaH3AwZ9o4tywi
raoQqNTlZqp+b8wtoN+0l/49sulqS2aKlMZyrZKbjcOVh9VlGPYLfLVCArii61yy
iNmNE1xbp8sLZrnlymf/Rg0bFnsdb7seaYBgGNx0PkWPfU9lesrbmZwg/QBUi5r3
6J7EGfetZvLrRh7s1+ue/uJLzEDB90s6bn7LoN8lDX6/MJvxmkqxqo/wTp13XvcT
ubgWFtWznZLkOMOJqbaBMp/0wTQqu8TrkXexr27u91i7EQjbEdILE5sVHvS9CI4A
`protect END_PROTECTED
