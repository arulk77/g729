`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SfLniZhvIjH2dnkbUYNIM3zeBhGywufCkJDSchSEL9gH
uVQ90BRUWFBljS04dXesYORu1aamqYU1UjELCtLy0AzHnGwl9UOXIC14wAr/BO+t
NfGf+h77fvZoaeli5xiyBA6dqNEjQxjlXYMJphPFoL2mGbQ3nYB10xs+5DEoTbdp
7B7PjV/2/gXE3I7bfQXRrMsMrDeKGNZHHKKWvupBN9KkrAnMTTNfim0bMLg0vRAj
2slZF0frS4d93gsviCcFpwbzbdPH7EKasEuH8XyI+c35WPrsP7cBVfIxylaITra5
4M/JKKUGncTmzHPNMiX6mDhVaisKbpmb07x7Mb6yghfpblDwEgSk6BFF1yQn0S1r
gHDqe74RanyNR/zwOz5masqjwMi3XHMCST6NSY9vzxI/qGgC8B/BOZC0DhHqAw9M
vbRLrgxzOX/AyHnrQqhAEijaqUJ8XtB9++953T/YIxv0O406P4Q8Qt9Ijj+0aPd8
R+ZPnpSxe9RxWte70/uZF/3gSyScYcZMkX8i5dAptqCGIiCYnY+3IgCdU3V3/D4X
3jY/PphWWEueQWh9zcLmt5EzH7b4BEdwFThOBEkYqXtuCkWfum5L50wZaDuhTj/F
oMrUBuDzcZrCfQX6wQb7IX5/d8ZewQ3uH1aJq+cdtlCxbVpH4MRFYBQYf9zc6sAh
48lO8BvN2ummThcDwuGGyT1SGBuzRQDYVhr1/822yk+irXkytLiu1txFamxek9RD
Ompk+RXmQA5sG9lhVEuT+fGyCA+MHmT3TJ2VUSLM2fmeOBdCMK44H+CV9cLAngCc
Vl3McF4O7oQvhGa+MvXYgrofQfrP8bzV7KGyDtzEOgdCaYTeoRg/1mhRUCmw3igO
VZJ29hkPwnKophdWTKIYFebc37+5m56CB6gSTiMKYtxjTvKVNVK8rCejYniGAAcx
7dCLRcuNwA8z+YgtJTcRy3VihoQoZPWJKmYoa0ZIueAhdZuHI3DMqUha0b6AaPxp
PUUFuew7RZA17We28+b/czWEiEZ+u/xUMuVwdf0mQ/XvRHRPfXAYXHdzxShM1tfs
SKG3X76uJtVAOvrYrAGagk0HtQkqv9/JI2CyAqDoZWVgSfMPeTH9Uy0fGsAyRBLS
buLx9tX8vqpeHtBlVj8Jicn4vk9regpYU/tqPT9/HFfVkCnUMFIiUQxK4ki2+n6M
QWLzDgGkkaLm72wAKAIhSLUnHg8gL1iATWMTBQMmGWEiIlANhyQ4AaVG8jrWT/2R
cCVIAzCH6e4y+Vi0vGbKV8VJyXwAWg0wyxYomJnqu1/l/21tcmoHiJigfXax9OK1
Z6vJun3RGsYy4FbwDd7spa4o7uXO5EQoYVWgkiMbQ8gSgMqzKWcMXd7rKY5zJ32U
HUtdmz1KDMCSZP+1kVl7jokLXEHhF4IvWquKeXSdgEBXTDQJUSt6lJBV6rV5q7L/
bL//W6MK9X/8hDXr+JrXU1md4JI4qrkHX79ENFLqSuYHmaqir9kOFmT1QpYePwzW
UNUmroHppS/wkpvRtU5gbD+94ZXuq3vog815xLFwLPxJrNif7cz1WZpm5X0DPseW
QiSZ8XO9OhzQ9z7AAYSF8ocy9ewTKiktLwp9PvNVM3fsVMBmMJ4BEwEnDnxyf38E
YLqnWcfy3jdWqdY6ZhvH8ZLDG0QPxRrqa4HpsvE8V4nBoARecResh7Jn/LO07RPF
CCwOElyAuAWWeUzjDpDidlGOseWBiNMp0EMAN6FFsgYLq0J/RwSAsCX9jLYENP34
fQ1oM+RnJ1b3CNHRFGI6gk7lY47j0bIAMCnNx9hM3m0yEsShEnyR8F1H2bkcjB8/
3CLwf3UGYZTlLxNCr3qfuNF6B4+TCilhuEODBwvTNlaF5mBAHuE0g+aMajmK6+RU
Y4DSeSs2Sje9p+kaZqg5qX988acZqh8BvISb7u+6JwtQoobu3uOy5xHf0XcJT5/4
YjxL3hAMc2tufaD3AU9AO6yEL1myrlldB6glxi4TFlQoPHH18ebtsClVXc0hsdO7
6k7Fgpyg4PXNtlDcI/RXGN0HFj/LQN8kpD5Gz3SDCe8YSiFgdQWyb/H7xSjzMktn
oBptdES68zQbYMswmj8Wy7CoTGT8ubnrDYhW/YZGl+KHT7f+nLkfjc66YUafwdC6
RtUB/1C5dnE3oii3buKE6UY886i9B1urJHl3HN0xnwkKfb09Bvk62eqaMJnL+qkA
RKDYkw0EMuqcfn6K/tMLNJx0Zz67VEY5/1YqvxfOtECtYkm+gYZ9lMAfzCQ4lAL2
nZ4v13Tc+y+gXX4GtvM2/1rAkTlyIkNUSjEAOyaXhGakCGCHhwRyvCyZn2qlcOOy
RiIYSJFqn2BiuBfcEnse0vYkEbU+2fP/DIrPuvgo7asJY9F0iuKxil2mhY/ncLQh
oiN7/mTwb6uBOCbKS11tlRimCfbq17lZgqfCvBra7EqsXDCWcfaKnVqshV7BjaJO
eXczyxgomY0SlGa3xVe/5lxChW/01+80K01igCzfb530OwZZwfHRahWUxxUST8Ei
xtby2rLTBFFkyHPKos7YBRMYFi7S9ujOU5kbTg35RX816gOjWjBLXh/uoHP0i1L/
vXFSoscvjLIRjgJfc0K/Tk/ZNgZxJ92cVxb7rRmbACFq7X6ET1Sw4GaxzSF0nghV
GlhdN0ipKg7GnSVKs42vGg4Jdq4Dzbr5xwxn/vSbdYXMNGai4WGlGo/fMHGUtjRb
7IGz8KJzlndUR2uVMYyysZnXZ7dt4UXDK80mkUkMRn6dR/XC8hez/LQ4rzGJ1ade
+rJ9dGO4sF5scFOvNn96A+lB4VhM022hF2EQCPD/CmRYpAk7luOTKz46ut3HTdRl
/Zj7gxpM4d/xWTEsxSNpcZktCU+J4FuYO4oVOOGeF5Kw8cQeGJWUhTGpIB98+2gc
cH0uAEvHxPqwztaNb8iqkeADE0QTdgMJ7SO+wbgXeK7wjpHRmMpNr2Ep9p30W0IZ
VulKW4Jv9Jo1TSJobD53GVEJkNpSmlJMG0F+PYJ1c/Fpp3fjIBvQL5/WAF6LRMMT
PGWP1cl8bYASR423MVghswqLxF0pl3Gl5X/Iv2ipN78PjLSYDvUMNq2pXAqJpqmQ
za9G1/BBNW/XZkZqRlJ7hJ+DBUE3mcPE8OnJxBikqjvbz+grsmtSFQUZ5BLH4z9E
Cd6Nb7/Y4BAxF9zdiN8qCGuEX3FfP4spVE7tw9rs+DgmGudwYaMOlulhMuGp53WC
UNFsKK3ZfkjHnGMkpA/w1knLbS0Qx7fVcBqxXuU/m6LyNxxkCjUUBw51nmNSFIKD
eYezL87qrShh8R5Zazq4iCDKO0uMEkv9G+exe9nCpXXdlkcdeCxaAMcxK1TlBPms
9RbyJNHxXgcLtTXt8Rxqba6swhOHOu8N5IpuS9U+ofKpOOhxgl19pB7iSTGNL+q+
4H/QrNEyokqukIqVE/0X0kvEoUD1NiLwuS/qkD1yM1fBTiQHJuSWbkkqiFmRzO0b
UOztUtgLEm0X1SHtazgxTxzer0EEevFYuIeHnhwXUm3QR4jQyX3jxX4aM3+gapq9
eAbRTLpNFIO8XJUqbmAexmGB/1aLToSd+hHN7DDJp+R8T87V0zTmC7o2yUQiF0Or
BM2thJO+pYC4AwodiZwRZwlVmb6yekhHStEEzW3e4++3qJe28/M25InvVxM6rtPU
w3rUXPYikbjOY4MarkvMrBHfq2tXxT+muZ7Fnriwgr8ME1SncnIc/AW38zLNJt6T
2xKPltQhWpB5h5jLKisfr+oVGcS3aKbBEpZppO4HD1lbZzgAIp8peU1K2oeBk3Gu
An0fkRngAd9woxT0OhCwoWP+SwNqBxUK4b3prqq2/McraPTtDlYjJB2M0d+yP4h5
bTux2hqXwKo510GhOGOFE1soQSpMYD1XfT2re1bCiTJDeFvDmQxWtsMbHkQ3n440
UuwPFMveNNYGy95M8Nzku6yx96/0HYIqMIswfTTqzut0LTuShDJr5ZwR+iUTLY5E
EsHZQK4bP4U+f9FoHmu9rcm5vFN1aXzhYyx6tBgEx/S1kb6212MKI8SLdIhO0Pdt
lgKCOakGos+06su4cotKefwXiziocw41Y02MoCXoShvjoh2xOSHSNkGuIGrLB/J/
OlYvwNRAeDIQuP6S0a4GfnPprA0kkGQpg70JgZ5sy00GdaMdAHwWb9ME2vnBnBAm
MEoU0UrNRmlKFiby6xh/sBPIs/SJ2/gXFAAB3Y4yKN14hQIzYU7YfzXWMQHZTM8R
V/5rCt077ilCrt4UegBLS/WxyhBJa6+YOqSWbdO3UDsmEUK8+t2BCNyMKyJo9iUk
v7rbAW9gZeivdHFbjXmLZDX+hHtXaHvqKGUSHnpwKrLdmvNZqLU9HBSM3sx2fUhV
Dx1ffbWsGZzsYtf26JRQuOkPgt5wNgoUMRxdAFwETdpEuJpIUdnKvXz43DivbqWj
GW7IRykn6UVlPjXWA8IOOJ4eaNgfADIsCbXV0e2PuOw4ejMf/57+bCy/wC3IqZWu
CEv3zKEab1zWIktX4nmWqX/cNRNOwckCJCZmrkGKZHYBRuxmztBVgnhsyVH4eToZ
MHR9vN1Og/AmkewfRsH0+51WLwv9dQzOOXSlOvZUqKXWRuRPNFX+my1n7XUXl/YV
l5zpqt/fjbvZ6lbLTLcBfFK277QJWbkET8eL0+kIzmhz4gLhaJQ85SreyU4xNfpw
CodkmAiLM5XRKgDoqcKUBEuZbi1UESSg0+PJhiOnCO2nYeT+qOrqH4u4612IsL0c
A5iSXVsTo4M4YZpUE6cleMEUAgI7nfZc/eBRRBlHjRO7GWgtZgQ9e9k8yBXMlely
u5lA/+olVMGdyJ+hJP5iGXlXaDz4pbEwFDQZoBCCmMXVgYSMnulJj1KiOqPQbp0E
HMQ8HDQ6xuI6tniYd6HEeglmAYl3S7NEvSWjR4ZG9sHUZLL40HyS4MEnUjvp2UuW
ScGGN/sV0LqjFtv3cmAd7bhY70q2/zZLXKFEWb4Nkd+TKY1jBKLMpDYroWgPzoQt
XOwLPDZ4S/+qHWRRFPmJ++2LmDzLIV39BtXk6uxmk0y6NGJZb/UieZrdN0H3IBzW
gSCJx1260ZDzVEsm6Q7kUSTAaOBSQurIEOS8aFEJ+YOE2pUhpqZHq+Wpk008d0c6
Tst72JOnk2QowBwiKlMn/37wnyFg/fCrV7es4Kax/qrj0mSQjQT+Hf8isu0N8Sv2
11PlR/MR4Bo7s4qtubi7Sg2AwuzdSfiGwo47geO8rU5hdRCNZ33bRhdT0DibccqK
L9hHyCDauNpAEFGM2iJhMnRWpv+V6z/LXCqHsbenP8UPv4kTfXXBMYSop/gU4bNn
ZnjzZcibbYTrCHqdw0ov/1a3jFgscXUvPTN/bJJNHWkflWZSN6jBIkAxUVcAhLDT
l3WWkK7qQPSOpLBxEvxiNifNZ34glIMdgzH7KLd+cNTnON1VUQ6B0IszSZ0FuYHR
lgci0nkVrKRcCbUp40DkvA/3xuTRtbfmG816au3I9XhJ4TCy1xlj2B9sdntb5kyS
KCKAKTERSnn3EhrNkulPFNRSVCGDakvpRyaUJQIjO39MDgBvJwZ/ypmGW8vP+ZNT
T/ps33Cu9N4q4fSwGs8LJ/A6wqzzKSsMJNergnLWY/ClA6q88+dAb6vj4lWPFKur
U+UT9Lb+TfGvnKljS3rQ22GFUVv5vItJ7uEdEaakTubB2LmLKuFTV4N1vUEalyeF
Z+q+KxXxAPHe59RBRwuzpqrmUtIJDVhXG25tL3wLI/GeLb9MXVs0Ap7ryjqoY/gq
nGk+8rOf0n9ekIBdJ4rn+ka8Zohg30mrZ4QUPxlnO0fORHSNGNV8U8ySog+/sR3C
5qAr/OKqeqzRoks3RfrS64je9RyhJrgT2wFDdweuqk6o3kpimJv2rTMtIcZD/ggi
LyvsPP6lkplB/gARlSdlvfhjjzFfjh9yvwigovlqULyj1mKAbclAA79YezTQh6V9
`protect END_PROTECTED
