`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJjaJhgk4JmDvrxWngFBp3i2jtukyARdJuOg1Cv1MB9J
pCccxbVNJuLgOZ1ROE5JOxE6STSFkeBrtD7x5BUHaupLvviIZE2OMMh1ue87ukyL
XpBGUWdVEH6QnMsdraFMdrne2cb1WIwYJcOP0NUJSohLh29UhkC7KLS9U09g6RV2
HpW69fQ0v8iULd3zESB0yw==
`protect END_PROTECTED
