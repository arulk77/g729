`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHOa6td+WyxrU5vtdcAxyQupJebKpBZvwk+8UT1CPPTe
g7UWY6FY8WySaFquKd3HgNgeiKlBd5M7aCtK6ht4Ia7aJFVN2AOmHlS6nWg+021b
JT38ZY7phxpo6/Y8BkulTdaUJu5agF2RXAdzH9L7xPXucE/Lz8VNko1vE47J0U8p
dIzXuNJ4ZrfuRSTO1BiKLBpbxsBEiTn6Q2OEhbmTfvEI3xw+6hkRRx3wlH7Gvtc4
JpmKk/nyzSL+xwlSKU0F8g==
`protect END_PROTECTED
