`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QtKWwlinhP2kdAp/bUr4HyoLN/mkxcVHqFPFd8TQpRfOKzIb1jrUYv2/tpMYKXW
5mXDKYSvwqT2JBK6po6DOptTOQaQT85eAWd2JAOuHTXdJMS8cL4gwrHbiqtDzXM5
gfkuXLlT2zteu5ZwWhK4cGmkvoatcLA8/Fq0OxZc1cgsjghFimYBU/zNcU+SlLJ2
2W8+1iRhKxLB0YEMNxQ+mpb7jWhBiRBVwj3OOb9IUiFoIo3/VlJNwe82bxlzY5ND
N2cJJqzyDPk/fD/4W6qwLSk5Sh3Deal0iPasQnFgwQ4=
`protect END_PROTECTED
