`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiM2nRCPDLpZHW2IWaKarP8CQ2/PosyG7/jQnreDPhzGwb
U6dza2CivHjdplv65aABCxRaw2SECZha6lJK5vNXftwt35sMQp43Ery50WJhL/jt
xxJcel7Nx1gZFnQkvUfZknVMBTzhY6nT7Wnpy63DiEd3XqbmRVQ1jhSfU88WCNwh
zGcV6gRMqPfXIiARzzaxd4Vsj8ZQpXk+xd1y9oO/Gu7HF84SvoOSQfPhY/NR1yhO
`protect END_PROTECTED
