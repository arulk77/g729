`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44kzoR+Kpqv4B0yIMQUJcOagWlvOo949j2cWW5Eb3tn/
gH4H3spjgGdj5p4OqbA/4wzqYDJ0jadijKOCvnLTMsdZvKZHdO7DHfIPPeyQxG4j
/P4seyLpFx1xce6jYefjdowuAA04CSNdTOjzULrtsWRREOiNQ0rC53lOxy9T+qw1
ah4qhUNr9qQCKhCgd28C2oea59NRyiViQ4nE2CFjQGsD1SISdv/zgR68IL7XE4ZV
3435mniaHwdiduGDzSbafTG8nzi5myj5HgET+YyFBXWR1CrECUBE8Zru5Z6MUdmf
4LAyF45i7wGz00GR12izQ6wYFz4FhOt0nonMr2UXbCf+xiWeP/vHg2yg9SL+fvCD
jpCBsmFJRPuvQM7K7VET+gcZCzKpAyPZrXSEqvE/y7QjweD2UmVrQ37Of5Kn7tho
18iHt9vHqzOpvhRX2iewirPvo7YtLPJo6MDid0cD9fFOpixV3phuBFyuuK2RCNp4
yyJRcaaLcl9sL0kRPdm37OFeX1Spw7Yd/z9k4lejmLn9HqzvTo4GFY9YA28QSaZ8
mTVvw2aGRRi8af1gLeSQSYd9jgxhqcmXIzJQkVpyKStBzf4axRkm32uvR0iUOhsx
9/LCK0RMjKigGLBidF28d65Yotw73EC4UwtEfpVpgmJq/i05wzKRslpep6mTHc2o
`protect END_PROTECTED
