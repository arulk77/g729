`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEIklFotTcObyPpNlHacab4dK1jJ+nxTjR9iqMwQWGdP
bY/6rFfRaHxNwFxJbeIiDAqON8tprByv+ZgzJDai5dtH75EATpvt4gqqJN5AiONY
1nEV1Nq4An8Sy6IG9Q7q50hfwd2NzxS3cOAnkR7VCkSRmCotLXWwj/oGNFNOvOwV
hJwclLsa35nK3HJCHE5We8CGQhwMVtCEryH9ew+vc6Z1Mp++SfzHzvZ4v65isT3y
bEI+dV0RJ434F9tWUVUKHOErvVtxG1LGTxowu0no8JCLWd3yRocsWcxgXZpXyXOh
`protect END_PROTECTED
