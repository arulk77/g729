`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDPEpKvQAriN3adU6mOu6PHTJD+QB5WF5RRlkSM7jn3h
fXjicUBjhrL7aYqjwDznMf+qLKVeJYpATMA0qLRmBKPWMWLz++EDEhcHbQV+TNgg
fBTyvPTadn4RGi9bpVPDF1zjKdSIhhFEFunmQP+isxGHRpEM9Me2aOfLzSzEVW5G
CK8a1f25hOxE8Dl71CLj+34tEVmk7RYlDGYvHw70oUzRY9pu+6E+HRty7liYEQjH
w74fUC4EqdoPJZEa2nk2EkhNRofmrkETg+gFM49+UMA2zhJ+RFg6PfBqX+8gkCuB
Sizhah1ECVGIYOoNEdxqbKVLplADDvpo6u+0GYmqwrFJIAR2fTs6lbLl0K/aPxng
N5w+GeQ/8RSOejq+dAic5uew4560MIU7BCJCPiNiIEZvmC3AtAt90tV4qq4uSQA7
lsJ7PWLPyxx47Je5vU70vzUGiuoTxSzg8hvOFkqvb7l5tW2gZ5W0HpAb0H5p09p3
FhXtDBA1vGgZaGaN11AVEBmWYPwAgwut5ZQ1aK1pfg0JrqlFdSH8oI5/BQFK0QNF
/2aNL68z4FUK3GkeFC8WIfHyxgzm5n57Wnty/X7DBH8E4zASlZ8D0zatJS3sUfTN
cjj+tcxddaqQG0MFe07z8PDqmIrOSdJTcNWuBx3E8w0//QTnOilsRFUKXSn9i9tn
vxdTmk0eY9JlERQsX3U/FjsvgJiGPTemScsvqCvu3R+qqO2puFDT6twY2W/JvpwB
DcGJFNvh3s8bvN7s2qPk1+LltQc7nN5M9q8g5eOUUj50xGmlSKS0bE4JML2X17y1
B9RFRq3/EBiKDhRcqR2WQ0qYyRhNB+bEnQje+WSwDt4=
`protect END_PROTECTED
