`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEhAC7OLGyIhO8bzrAy/Sv4jzZcpuwFT2PjiUWlf9VZ3
HpiAZofYmDZdLeNYHIWdvITQ6AWLJAd8rf4DA+LbNPzKxgWDfYC0fjLHCez9voeD
dEq9Hc6qJG3IEnhdohGnMGSIf3xClx2YlukgKcmemH83zsMmTUCC7lX2ZZJ911yE
HvfRII/DTtv/ySUJhtgFL3HFiiFt1VYsHFnMwSauKxlh3njLm8DS32M/RCVVQj7y
Y0d0n6BhOMovcRgsadrYfJ9GFwv4MqhpX75xHZbj1sMhWANu+3/+1BG6awaU9Ymo
1TaoirQ+aziPIGZj9z/vg/fQ0mkVL8uH3x8AV5jj8uAUtZa3h4fv/p9PEbnE5dHE
2KlkuvlzydV02F2ztNUQ5tQt7Pk1pcf3YeZo/PX9rZOq/AlHhAEJAEgV6YqHmZja
0pGM5VF+Oip9bIixtCaMqb6AXl7c82FvGI5H98DRoZb8CoVTSQVFaLw/5dxFKXSy
jGNFXbIvzffvzdkKvUe8pQ==
`protect END_PROTECTED
