`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zNffhWhuTe4On7QLmNxmA10wYfr/N56QFaVIwomaINe
MQxF9b091s/5GlVNUh282AzHAOQnrisYpm24Pa4tJUIu3SIxMK8yExdpJ50eGYk+
0l+HeqTBrgjHudcc+azPIWe+Eifr6zBAyw5HIR5UUO+LcQ5jz3uvc3r+C0d0fSCv
Or91iM0xC0Io8CPKxeLLf4aBinOiE+iysyGbS+8D1os=
`protect END_PROTECTED
