`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48N0WIPWV7Cm01l47b8RUrKOG0mpAfbp6XTteZsGsKe7
RJXQy0zK7rLTLVMH0r6N3O0hVWmra7Ptakj2SVRo7FWg+rQZ1XlCvKUFiTmTkbOu
/3m0XWuGKhrzOCy6EabgdiuCvD5G2njAw3JZyR2X5h83QibSAjOYNAHLQERJJ3C7
ddD9tg1fOwoNSmsAK4gbtmEUZNgbYO2MpFVUZENt3C14e07KhWJBY0BWsOqorOKC
6jeSG9SxQLgGzmTHQWBQDfrvxIBT9SZjNEK2IaSzf2otboxXW47hLIvju/CMa7BI
6SruZnzD6jFrc19JnHNkS7Zp1jTBdmQdEup4RtbR9ruJaZMTP0gARP9Bj3MvjJgg
WUzx0XTEpErKGVYR9lWp4A==
`protect END_PROTECTED
