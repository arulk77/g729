`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePDaet7lwGzFufRRp0Va1lDlE1BVG3dndHgZAUrmZT2U
5kGq2V7f9Fc1XxFUcDefx95/qY90Qu+yNkiPWkIZGOwUKbtQjJ9D3WU4P5M0uzJd
vcFGKCyvF3HUfNEG2eT6yJZ0zMl5VPNHFa++4sFhNY5qOhY+PP02x+FU9I+/2wTN
jl98E4tE5tgOjwk9cRn6bxWibVankfVYThsA9H32VkS75vm+SXqSc+9mZg8URzjT
VjC8nzrZVlZwb2hOBQYTbxUmOHvX2HE0bBqQtQVQHx6fr/ikEZTJ6mi0bx9PI3lZ
2RMyIg3c1hxu/ovJdmg9p2N9wwEnP3nk6KclwIa3nZ8qStDuBKHkhCTexqHsJ4uc
A1ofngbsgBp/MLuM4QG6792qYBMGb2MCAG2vMWrnRAptxVaCMR79ITV2p539NzNL
/OqR9t9m1sJK34y6z2K7RDGk+y3h84hV+57YOULfiNz0ZYHPd2ll+brgpehD+lsd
dVzD/Cf5X/tEj2kc1o65BaUGHx60I4d2U6hW2/PWxvChsJS4CbEWv/CMTldOSKTd
rmLHH9lIkoSsq+b3kCfp/VSiWNBrqK4vGBcBd/3Q3LMHtN0wGY2BrEdUB1YNnHX1
DGi1rzovnqAOqZ/xRXrQzglJGaRUJbbbzEhVpmfXYke1kTZyCgFS1mU4OrHqq9mm
/pHo24bB3/RC1MHuw5h3i4S+HUKEXdI0BAdWOw63SU++qsNNLB0+TLxU6XLdMLsQ
u2zpiFIsTzOiNvpXKJcqxPTcGhW+A1yhYBynrLOmc6/5q7Yj8rdk3Og+HOO2aMlP
5BMDLa8Hw0fOOfxekGubtolmWQrY3rv4w9+ceYfWKYuoOo23YYkrwb81dg8bERlg
y32f319RUT9VtJjgZl6eaGsjjlPBB7VAxEZy60RZN8GWLSJhhEdAfe507Jxuy8Pq
th/Q5PtcLo0NfroIOScHLgmIOsgvo+7xuS5XoCK1OWVh53XV8iz1bA2PwUnl0etq
cPX/a1SZImbcM5Ef6Dz6F/k4DmmFAY5JoYTROLb0JbpVppRp+Pl85BoDGRqM19Hp
/AXKDRCd+QSfqL7RAAcFl+xuGxnOnaztDtmafTI5Z7Dr5FIoLvCrSI7Lq0RrnO9n
+DbI4r8M2WDoHv3DhZ0KBvlY9asoQbJM9kqqhQrsRD2biWBV431LsMbcSENTGdHG
87v6nD+1lvzRk85JnjGs/wTA9ZF+TWoJPDjQzOz0h7h2y7BdVr3CZpRteVQbq/5k
yUz7u49/Pn5xS7Bq48H9kmL0/Z0FXVr6Di1qwDpJ9y1+qQ5PR9R6BKOwkO4btN5x
8cZYo4TOK44EIWxnZ5hwV8JLWViGqzWU7a7j12hJgKCs8STIIAUh2xNx5yrlA6T3
Hvcmb5V748JRJsEyTMV1+pnILSj1aOb1H/svssCFntJq5zNJI6wCVvBH4BgShjik
/brOfCzIx7DyzM2XCiNPhPjNFbky02BMeEKXHfjdva3F7q3bjU8qT5F0UbFDCx6Q
u1GvB2JsRyz1RPD9hnOEn5t0qS8RRCa0+mO2h0gI04KdxmvxFyfFdpC0A/leS2vh
rioYDsc6gjr26vyvDFslK089tVZ/xeIpuitBpqGPXgnoQytKrk5v9Xdg6WRTBezX
gSixfOdR89ssKYKASIJOj5DkzoCFm3GTiuCDyz/5V2Ic6G3nRjO1W2qMXEuqKFKe
`protect END_PROTECTED
