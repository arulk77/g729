`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIiyaqvgK1FgVWz4lFN1yTiPXrmfKqaD/w3hmEi5/Oh7
iX74nqknEj9tOvtfGK2d/NfkgQONI/0lKihrUJcql7w0r5lu/EBJ6OPZdB1mfRnm
VE5vPOdOOeMHedjtoUa1Xaa9pujro+5e+SsAXWllwS6HH9cf/ICTOBXjCccscdDf
0ZH88Pha9KbVppJHOPDuhs2n+XMSNNzvicAkQ50GZEWLsKlxwTku3EJ7B2cCAJH0
Oe23nZkWaWqSfCaxfOKuAK7YeBXoq2iizg98SrgmDnQ2aiMI9NVKPvrCrLBaFI6b
+395ob/sBhSez/b1C97xg1gpjy2RniYsyxofkQt3pe9vVFLM/G3z8Wy1tlIDnZMK
XChRzjlFIdvT4Nfg7zXJy5Qnfvwaf9ZH1+OQ+IRyG7Wn7n75AqpEL9xbcUbBsc4Y
jAM/QH50B1UyNrnkJTiM8RvMBxuwFvlgRckusCTdCOPFZPyQ/w27hYAk8MoUgE7o
`protect END_PROTECTED
