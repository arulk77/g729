`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCbcRdGLdpJ+4BtcK9upK1QJUskl7p4NpnNtOxNwu/Lb
JMWZ2eYTSq0m/QjMrAPEYnoMHeHfqsrpFkPyqeL/ocvguI0DZILgj/eBZ/mj7B/y
/H9Eg6iOaEnZENuYvVzeZlEcgtiZLzt/NvwN7rYxml1f3zEgLuq1CQ9CofsaeLXm
`protect END_PROTECTED
