`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dE4T4qkB6lkHZHoineJ3tCA9n8GqowM4Cd5T3WgDGw/PiaZod9zPJknXWTaX5Jx7
Qj98ymSE2QGobew5j1EwgXutQqjX3ZeJS307tx5uXc90ZYrnIp1pqhyG25i3hR4Q
`protect END_PROTECTED
