`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MnX+Nx7QrY89NoEYER0MGXXsZLN9I4IYLLAAfbZcjK2J5znQlpji5pLjhnOk3jvh
MD6vH7CkZC/G1s7UJmMTTJ0mG8yuXGkmsOHKoeD1s1FyU9SYWQzsLPNkVLpm0HGD
evnL0cs9A48pdkIGmlCR+HlgM2vUrlKdshNCObhlMMzvo4cfRRTujnw8RpVrxJTq
bJTu4MnLU7lDYkQlrgMYCv0wMaR+4IPtKAyJzl1zO/4TWz4OWk+K7YLFR41S1t5v
Oy/cgcG6u4h/Ez7FYZ1QYB6g/3uyrwBxDM580rmgPRs1VNIXAS/eLAPik99BPOPn
78vfd6csEUdpC5dFJh4gD1B1gbjW+ZDpqguinHnKvpsENJqow0pJ85qXRQVp/H78
VY8GzxACMDzqdKi5paYNjgRlT/xEJKJK2qtiC3XC2WGZxVf2Qww9AheV2EhdPz+/
thmgH9VX2m5e5BlIvuFmCt4BciHgTozM4ziXWAigzh6pIAFwipMrk2TYy0TU+G07
8KtbEqxfadwhUjdOGlv8O9bRekaWOT1YaGzvvxKAwArPyVY8Tsp/QUtok+Mh5yEd
GtWVZJJ13r/AWkfG/ubJJXi6KjBIpnGM9ZtzvUoXq1bKZvg7yjcv7D/m00c6Lf5j
9pZ4muZ+CrH/Yxa+mKUpttA2MpdHI/cy4WZf/qR5JwXK42AIVPoGjhlLnYSCcM65
GGQ6AgJrWE7XszCJ+ZzaIkcsozp6M570wpb5EsPh2jrQQGKdYPgs6ELNvGOX9qO6
`protect END_PROTECTED
