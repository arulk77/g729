`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePrJrX+WOMEJnZDvJt9qzQ2rbBmXUMNtJNj/U6O4prMv
CT9lwo80qr1csehnVX7tnldRlBKRri0Qa8nFbzt91m41M7cEuXR0b43ph4aeBKEu
DC305ZeEnHHOfM3Kj8cynDHTap4S8XBlc72ZYLGiI4tviV73Ud3vksLOiBXDR4c4
d6XdJMY7P/FQvXGyCLUR4KFU9YBsT0xRRtuX7poKJIonXf5a8mZ5PSHP9iiBPBdM
`protect END_PROTECTED
