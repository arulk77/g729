`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEqeHpISNmV0LBvJDl3VA/hEFJ5y67ze5Nvpfknqx8t/
fXeNDBJ9Yzj++L4AUwRzX3hpvI1M9Inv0qVoibJ2XGYZRmNjRwP3ODPhVchTrYd8
1G6QKqPWijdERBBW1KGDaBXBf8i4MsOfPcJpc7MBHPrgPglCLYgwn5OHcv4ZYRtH
xyxKSe/Vi39eY+RiL5jfOZZDN0JEJaBq83NnlAYRCvvkxzmVpKnW0R49xnPbJAei
`protect END_PROTECTED
