`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5nipKXlauS5X6wpsjRbptM8J9cIQrzS75i+KM0ihQ1pW8Jk8sDaTh75rTCahYiAc
9S5FSiURskPtOIJ6nv6vfH/kXp7ib+KQz0/OGxg9kZgdZBWGenzM7QeTv8N4gF1+
ePcn2tz4k9Yhh7REOiZvSm/f9E9KGDQOU4K1w59IgRTyvNlfXPLPm5DG6TyH7Y8a
IwW7YVb+WcETTMKi/BaFecX7RjunM9nhC7QHuePqQByZTHqzjW/ijZvzjA9wS4Xp
osv/qez7rRDY6/NKzum/GJD/SOSp2DAEclnd1P+rKQXGWeM2hFjBfhvsL2MgdK6T
wZswHB8FVlTpLmf6gLu6y4NThcht0v8GPjBCM2fQ7JXcJzGKb3ai6jPYV39BhHQQ
zKHy3J/7t9nKrjqm48BwwW+qGsYgWk9ghYDypTwgabTzVRKjuDjNUAb2l/w+BxIW
kWJJoIsQbk9pF/4+/v/qflF8hrb/7RfFD9AMpC35DdVudj1mTb9MuTTnAd1yZJLE
FDFGtCBd8tHGnM/BXzcxoQ==
`protect END_PROTECTED
