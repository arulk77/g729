`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C4wE3OXzJkGR2ymih4jZkpxC0U4g0v5EWeqr5kr9P83f
EP6HtBX0q/e+6scvZcWgniQb9jVIsFJ1M5k7emMMLvf3nkag58DojLsJOQ8CBkds
95W/YU+1NG1b91YrusTQUjmVLYSAWUySADtfuBq9Q8x6MYAeDvQZzpRPo7eEAw8H
EwmkzGA7Qa26v7d3wHXgOBz8aS301RmIwYTZ42FMe09795xY6Amlf5ughnRrMaWD
h3S+YBHVyjYd0l24DzJqftfoQCHmL8weZ4ZVEjJfWMr4pH33M8p65nuDIz6hKz+6
/xM0+rvweienBcUnTeBPb4V6/8j7IK7jDFl2lzbvIuLOj0HXYglV8bWCMZUjiac3
m34vMDNL4w+rVwEibqVK+JhQUfcVDN6nEop7jtNXkQ1FJfeFByoMHU5tQ7Fojw11
9Xcibb6ShXGQzxCyzuJlSwiM6We7W3XxZ/KyeHFlnJWYvJA+zmOQkKp0THcpw0YR
hviE20X92e4ZozDTNHQkHaaCNN/2ZeE2Awx5FdbyLPw=
`protect END_PROTECTED
