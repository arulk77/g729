`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YBw+kQ02fdUHsoUcoYlZvaRLKZ5FRsuJMJTtHdDXUBCC5vCHHNidAilbwxwWOyvl
TsK5kqrBfHdoyyVSFsGy9DvfIMrpIRjnOyAhfEBnMVctm9VVWTsUQjCr/Z+kJOEc
TiwxJ4eF0QxtWMapoH215JkhtiNwc2H9k3TF66IZ6FG40aY4L7v4RHOEy1NohkTC
x70mIV9zrVzQYl2+KNB1ks9gmB+EJkCSgZTfwMTYVtSNjXdGG2Qy048Uc9aBxy6H
zX74QtyqYca+g2CrlfTbj+8Amx/BpNytWRifzlpAqstc5AFYD1OVrIiZX4otk8Qd
e0RgBnoPNzOgv6MCYwQzZoYnZyAGeqZpzCQwBKLQr3Q=
`protect END_PROTECTED
