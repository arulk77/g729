`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Sc7ve6Tgjwtdfb0UXL0VwJvzBsIeSTcMtecTNNfQAolA
jXhAFmT3GTpTmLhdTc+s5Ca3Qb/Qx6loyAw5P9Fo8XYT2UWkpoDqhKuj9ul9LprP
jmlF9tEF0tVql+OWWnEnOkgrfqti9xwmr2wWiddELHQlogXDGM3GCPeR+Fw6P/td
E12DjycvX25wbz5CFO3hzE4fvJjgBqVCi6k3h9YbbmN2izQXeh9wtP5rxeChKArL
YX4TCJu1uvkfMbz6rNA6gwCzPdqWkY+vI8Eh6b/IxTtyzGl+2VTRJzTvxXXk4+SK
FuxI0k73Ofko8cTbdZpD5nw+Ev5loqIbUvZUBi5xhq2vmw3Su8oEDtuviPufgHvk
WLgtMPWpq4mcmefa8p8PY77JQsv4WLhLNdxKc9dDtzdvP0j/JMtpQdyzX0ROPQBn
fSWOtQjF2OqkDTj+NzV6KHXg91zY9vGIR/d5Kguds+kL4mOWUVXzzA8F0ctdbX24
knHNgqgouFuO4h4Ytl0QMhC/xXFAgjJS3jC2YKaUhBLkZDdIWMLGmYNghkSS0kju
YsT49YkVPeSd3EfX8t4xWJk5mzQQnuPwiRQs6IqliWI0sFcOcdyI7XMzJDQG1Y6Z
jQGCO8pvdimzeBf9YYFpCa/eJkjn6LfMWkPI7oP4f9TDRQDbohQP2ocJe+rPj5TR
KBxjPKq41iMYg1EgG0dyS8opopZUL91w77C1cB/F5YhPPgiA/rvs3hH77kLHD+Ym
`protect END_PROTECTED
