`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDkCbHrULIVYPTSL+y06HJDlkWZQyZMTQGOcV6O/Lca/
ihdIWa5f7SSzJC8psJ65Tim0K40pVq2kFDbMkcLrPJdCP62k0s9F7kP7wKVZjLV+
J+oTQs0IiRX5G87wEm3Uz9/igMgiBWEgG/6w5mNHSE3A0vgBCQryeczgqEeK655x
MMRWedvusDot56STFltmlUllQ+3P63R36zajoj4FYUUQKeh6RqM+crj8wi+J3Voy
`protect END_PROTECTED
