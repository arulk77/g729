`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wphN+/j41rqxZomFLoj0MT6HROuhwh3QcoRxZepjk4t
siaISDkpDRKtS4KAe0zrXuGllXPRZ0Yf86ZOW08pwg17WPOOVGMUAJvr1nMevqk+
K62V6o5RRPhh3DxwNGUV1tg7tAqq1PJuiyDoh0b3in1kv4T1UYiY/u3H1VKRr6oh
WJ/2oowazsnOSdi8cNoAKTIceJi4gljM//V8lzA67248jPQ+6gTWhfaxy3Gw6Czf
ZXd8aLPKa0bmOuUqUi+oqIUT+HzzkEjRf3J3JJgRiT9asX9j7OvLEeotFzxO5A8h
qokjrxIEetphEEOeF4KrXw2sf1+OkG516SSvut0VsggXkVoK35LPT2UJfLdSUwNz
rjzm+ZwVsnn99aXcaZZ/sA==
`protect END_PROTECTED
