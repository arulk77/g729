`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C1e297i7a/Hz+F/a/9REMvPEFsFdanAJk8QEEhhXkLW1
Y+vzj4CpfWYiHHFTnDCEZC44wOTcDDj9twTiZ59ldWnUWPxxTsbzzDuVffImlHP3
L/gig2GIDVvafGCwRjQwGkTS1WWB9HyJPGMHcxp9w4vbAGPztncvWquMUPWN78bX
q+3jVcXPC3ub7l/ukDBsgynIswKh0FPTaPekOuhXDrx6JLpzWQhlrdzYtY8z5cK5
`protect END_PROTECTED
