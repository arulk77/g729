`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wgsUaP7RImrwkdFOOECpXBBvxZn00LxIOKaQgBliJn3
QdN8OwwbWxkOIIVOxpmBhskqjl3nj6a3PBEss5NTGX/fbY5T+er6MDo/EDz1B1IN
lyZSkFs2WS2a53ug9+MotpEoFLRTJYNd8DlWAon8RE65oqHVLB7lTFre5jHHUtIv
7t8N25aG7BPu6m0spW9NlA5r4VKEsNeBcWHohi5c0TdJkXGzLo34K7+ND0h2qkmJ
piJCUNV6Qaf5RsrsMKtAjpoAi/GPPJxTZK5DAbgz/+NT5kU/UADAdtMmLjumW5De
n0BgKkzxbbPlRvsl5LFEZg==
`protect END_PROTECTED
