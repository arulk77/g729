`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGuOR7rO/DCSnM1N4Sx2boL/Y3OJ6BO+eJJyTJhbY+JJ
fnk7+Va3oroIOc1i6q3fMz5XzWGaCUGNlRQKCSLiggniiOCS4Qo2IXiuKQ2UK6JW
LCV3wGMS3ldjKF9CDOXEQTvxyIlCMC4bys8FD/kcljwoEXE3X5tHhkfqpkDbbvQk
Tpg7UpNIIYLfqg07B2zroNTWJDjILjekjkRMBOwJ8N59J+UGb6yju9JY9SOzdCtU
+ca/QRGEIlIpe+ikRa1khx4N1LRCpoIx+FshBApZjV6mydc1f/iPLUWEoC9MvJt5
qEdI5pubNFjMF+aoeFtIsXN/9JEPwwSCX3mmCUICXHVKWG6L7muhfhvVcey//A6X
`protect END_PROTECTED
