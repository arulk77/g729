`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49xhcwYy283uPAD8kYmJ5qldzBnSju4+F2KyVu9yA0cU
D8NDvL9mXjNrVRk/Pzsf03xL6Yf7BudWAtD2Mi+WGy543vioV4QNFQNgp2cBQ/8J
tdANug1clBoHS4i1WMIAHQDoFippwV3NCPdkSlFKTvLKsuaRn3HeB+WVYZ04UNTD
HgBEasnTsYWBagZ9LPBtkm4E55VAOriia7Oxotx2VLmBkTPP7H5SChCTtHZLe2O1
dfY5o5xLW65mMFZ/axVXJDIenwPMGNdR9utK72EgBXpoQyBzy73WJenbYzoaiLR1
BBjfrBHW6rL600y/imbSD54xhWPWjBkJwDgxR+bEA8LETt8yRky2/N48OgmV7GJ3
0jWuvCG+ESoLxkBk0EY76Q==
`protect END_PROTECTED
