`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ1HBkkDqtiDxgHT8/gLsgh3dYLCyo3PH1rOZh7zUItv
i4TqpTo+Qg3OgYBqoPhDdnesjoIArutdtitIQHrzbGYxYcDBcWOJ/aevZ3v7ywkp
S332e5XKnOY4pdTEWqnp4L0rQH37pTVTcTEFzVQ9YiKlM1OiTfMzhKw1cnpd0YvL
cD0zyeJm4bj0l2xnAYjhMr/dxMOZ9HXnYGV6lbmlvQfz8aLOFW8IdY8ER+xoX8EX
xeMtNj7oxVur+6jrfaXsi5EB3RXc1yod82wKBnJoedV4zOn0jgKCee3q3vMd2Vjq
dslwB3F83Z1xTKrrx39Q7Bd/tYE2FWUlMxnytGHBiWyZzAMSI7ikfT7CE6RdboVY
WlRSMdxh2Oh+rWpgwJ3cq9jaWkQb5oBgLtiTiuF0qmlGTAwZcnrHtE4ghEqkpZl0
gKyTu3fF397On6CiDvslCYzmLZGpJRitLfZoIvl6aU2Nt5F3DSSuGYFgdduBIGxk
RW0/l7QmdtT0FNJY7wAOkWuyqBn54XE2fG5hykpOhvX+caeqclVmidhY5CsMqVPc
`protect END_PROTECTED
