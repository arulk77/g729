`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHAYqbVyDPxf2KN1yYSlyMGDyzCP1oRejb2huyLYt8GI
tTmR8wzlzbIUaGbvvHIbxaB78B0IKV3vOKNgDQYYkXfmTPUui7WfHFxoPqn12sH/
HCwK6xIfuROP5yLckOgRwj4b+Kng5jyAFQ8C3VkX61V8Dq/CNsxDM0YGUb0nOn1N
klB3vP2Okxk61As6czwTsCkqiChA4mty93inYV0AEoIFiHAUj0g8vNLzYpb+pAKU
UVcCOFdJnVK8CvUTQwQrEOdv8uoih4xta/nq7JQHqgKKcVNdLtMr5zWj8+5XWckf
4/Pp3diHkYRy7kr7aMIF3wmUn0k6swsz4Fi1ABDQ8+s5WhAiCVwIvzsXK+gNXW7H
AOe8WZzhVcNXCS4V7BdIkVZgCXeXq6KVKqDX0KM2WoWfatXm2+pPI7QHLNatkp/h
ihemyOEhrhppq3+6NWRZbL3GRECS0OoMWr2emELQUOz7Ex5A6G2KfxdIPwFOG39I
`protect END_PROTECTED
