`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMkn1pzEhCuolAeoAcchwV1LhxHn2LO/DWL8aO/rLagK
8/USEQAl4qpUI9ajUH/POE6Pr+TSsX8gEYkQtdhTVjwedrw9wL6wFqji7EWddiex
2Lr8TfSsB7mDsxICSefrPfzNAfbCtHmvzPwrCdY1Bm77B63EF3Mj/biYCII/Ax4K
2Z51Vhy4v8haYAQOENnxOZ3t2PKLdcd6IEzO2m2vhv89sa5eP6hRBpdkz0YvYMHD
IuGyQs7LifE65XBv4IWtZOHhA5JWvW8vfc3hmNK2Eg2mgBcBT6dMUdKpfWReCfhz
g1C+cyotVpIfo+yyZifTbD9pGrOfr6RvpYgaZzoeoW18wJ5pN40VlnhqJWnPVzQL
`protect END_PROTECTED
