`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SdU3LzEz2PESk1vqUeJquDah0ysvlRSYPOm3s7GiFBsv
ixj5gJ4WqjijsJWhxXr93mKGQOo/KesTX3nSFX4dtRg5UNWXB7m1ejHYO+mWWt8m
0PTqvU7Wv7ZjbyRgX45eB+fRTj0nyxBuMXKe/GUmC72r3aPRSZlOM7t8Y7UUh2Jr
QpL5kTiZ6cZdy/vBC3loHPmCoarxJqy429L37utGJ+SfuAchHpb1k8EkctD6NLDu
ZGjr1GDWGVeWqheHJLD3Pye0IccVj30B6dtYsBcE3F+TJpXTve5GbPzlPocTrAeM
JPVX1Vt6s0A8F7XHzDmF+xKzWmhrBCC8320sYgcSPinc6ZUw1MQSOA0GpjBUAdLN
63oRgypB57v0ScRNcRyDj48fPsCpzHFctr7gt7Y5xxEJ21Fs2YWCADQuq1fKreMq
ASfV+f6jcmJIV5Yr1Ak/8faG1P2K7cbZGnzzkH43IHuAiZiLD/HezYf5prWGN2XN
spUv2j7ILuI848hobNZwJjvid9hFVTxucSp/N9XYqA46ZjWuxb2RyCxeiLS83VUR
NWn+dgiOIamLFhGlyt03ADTQJBgSN7FAl6lGXWXjJEEVWHAcVhQlKqaAjJfBYDdA
dVLhlA92SUmR4ayk1yN7+DcJv7ecRQ0L+MGFhRegK6qGfLM0mAZ2zX373wI3PGRu
CmcmMkrKaH3URgJRfGoom6xp5wrf0L1OH27UWiIf5FULbHRR43C+LOigVH7HH/WJ
3nNA2m3M9c/4XNiDbxoHCsNOeorKXvNWrfqR4HnQv7CRzGhWgEGh1vhXniIsPy2U
T89m5uekg3u+vhHW+/3wUgHKdR0yRPDsIpcFnF0sBwWnpPt6EpUNrgd+wXB0ZaOF
qMr7G7/lV83TOW31AZi88g==
`protect END_PROTECTED
