`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3Up5RRJnyk1pd6qrs1+KcP9gg3aSWzUzBx2KYTrI58A
CzKXBPTYi9xbnVvRKSUNaphzP5A4xhw1pAt837zhEsxY9JJve0LCgYXZ1hlcC48S
SzFgnISFClh2bKKac0sq+dwODU7+wuvCfmXU+KFvylbwZHOYyEhbMCo8OUzUtXpH
zCgc1HawHQU7W/QfvmblJnXkcicjzfReaQlNcMw6KnWWcPx07Gfdyb3AhBiWIYz4
dTm5cs3nIF1bF78P+hX/OBFgAlabyx8omtaJLTyNiV8YdVeFv9/AJw/UlEWXE/rO
kslCrQyUEzyxvefNniIbDi0nr3dB25lPgt/jG5Q7dBypxzN9zU/xmbv+OBx8++Mu
iM547qZyF0IxPHXUCpKHxyQXaTO9XYUokfrN1iIPdEj1X0VjSFLk1pwh1SMFR5fI
qvdnfEb1FmX6grEZmtjWKLFDVeQh3Z2XvuqUzuj+hblvlQ8MAFfRG8hp545eQiNJ
qNJwhXDozuc+kqpEIleAziFDZ6pZXnBbaj70K2z8IX5V3C22u8dWI5ra7ek+0+XI
NGpyNJidMIb1endhB60/wzDxgxmTJHDRDQGrc6BfW6U9zkr5CDGUYdPWe5bdUPtV
sE/MDrbPNg2PiLBz4D1jC7ZINY6GtXcg+uvrvBmDSu6H0lOZ27zfZTXO1lEY+TXx
5ZyR7XlpQHI1wLkSD0fJy8SYQAU0J9/TCPFh+5ChQAn1P6aCgaiNW9FQqq0XwOuP
VDVqWlKLC0YwzUJYrdrAWSm+aYAJS8p7L9l/+j/g5FzrHBJAIB35gZnNbHJ/Vdij
cXU1AKO3QSzbSYxKhKnqcRTeC9FPCYqNStstB4nIGk2OFDN8QZkpezYG+KGQU9s5
5q9OUU8km8o+lRWh3BU57BYuqEp1o8Ho2NbHT7d04dXl4u5bXIwd5qnYnuwK2xzn
hb+Qq7nvPHG/XRq5/7kGrlnNfYD7xvyXVDbbcQE6CXzA2g+925crkJAhs+qaQO0B
G7wHb3Y+D5oQMjxjV6StZIvE6Dt4SzuQWK12EuJ6RiP9riiPi+tQ+tZruZUTwbnh
ORMsf6oiE749Ih05F1xf3Wu4+iWCeZqFgvV4DdP6Ks69HKlwxXXgDVQV9C+mzxM8
TaIt6QRqwsOipbNC2YzccGYXG5nRj75Rz1DBQd2tPrnwWFGImdzwTN6z8Y6zSz7J
wUu0D9u+hF++g7ekLJykLEIoRwlTqvfSkYeZUmH+xshCMj8fsremYsRTfOAyMDiA
vHmupXR+O9xzZdkA5vvUCXUPuIG7RcXEF/E4/zReb8ZIYat+ZYrxjvt9Xflv/D9+
muSTihREDuM6tKtr3a9zxWx+F9nUZbY3/ieXi1xE3wnuFyfyPjMqQeApyAeHbN0T
7UMO0ZMrZnFl/mdki4vWUpr7CWUF1JR6Kde2K+DmkMSaJzkIOomMLiMd2dRgwdl9
qGxSQX4117GPDCM3Rexg/UE1xAeZv49+Ob1kTDCw9o0skiDyqCs5Ikckcik5wY/5
H+be3UdrGbwI2YGOrVN6rpRnV2m1S+d9vkpj/HLkGWzBc85NccOGmRM9G7+syMNa
FWbSQdOUfFdTSyQd06s6F0aW7X/++bDzbD1xNWUfmIelbhyN4LgYK1rqVJiKUVrf
4SjrTvLXzRtft8Xa/NkAPYqyWEMqBKVc15TZTTre7PBgiRplvjUHjS8mAp9tswo+
B3u4715miBTRuIN8l13E0UOcweO4fuWuLODkrOrf/SUFueFqAIV4Bo85a/YLYTMZ
Hla8lNTkTgfOFUvHYO4QBixPZqpXfv+K3AqZT8j/P+EUplnUru7lOigz6RHUis1t
PhwbPEYeNUZx5+OSUAhNoL5ZN/6Ru3j+sr4bPobQGONgIKg0fConBLhCPHTpJhom
5cMHLv8Kquftpz8Hfoxqa6gnGxJHoR7an8cNpor1DcTMnoqDurHUJatuSlA+asj8
VdbJwsAdeK3CRFk++zj89kvANMTKxGuYSTYlhHCIEllWa5NVS3tAC3OatnO9LfeE
oJcEMZ1GNfpSZTS3qUfGkFrtfJULeLqqTjMan7Z3w7r+rcj7DfQ1n8qY2k5Hs8mh
M2Z8scD1BTLEl47XO6beiX0eBdm8Nyxx+sEFTYROM795g0q+Cw6CN8FAAZE2JEjK
lD+S+0Cfi+9BhYirVSbbPayon7BqKFREfs8vKgLK97TFPfEOZ9VDzebvIYSO35gj
/Qn0cuTs5KV1lDedFbQdvVIVHjyNyjKvY7w8q6zaQLDUtSOgZeBCFJp3125FtHU7
mH2vXuGWY3LeoTlNl+sXbOkThv8Pbfj5pQm8Co2/lZsu7J9MM+MKAQW7YopACOgo
w2PAnFkMdCuHwkKtpfVp6qpw/UVnBHu44tILMzhSUukUFom+4onQy/gDBbOL5lF0
bM3E1W5p24JkXb6upOyU4nN1NVQEouCkpZvZptmHiKT1ml7CtcG88a+CoTFhFc6S
v4PYHOq3i9mu0la0Pr2miGdiCshhkDHvR+1GTS82vj2oasS+hi+vpJGHT4zSuE5h
/PF70XG2YeJMtfabOC/Jqv64i1hUuSrnUYWl3yuGXu9a7zE0AIW81bm4wBBUO/s3
myq0SQ9Tb2mJZUa3bnq85Puulm1Z0rpazm58tUwxuK5HywcwIoe1jiGH7LWI9Afc
RlOfxinCpjcdPiz80cthgIQ4cvmlB7OlvvpxuP0v0JbXlqBtYDJt5keC83qsbuLD
+33GmgXs8RPRX5krZipmIzadHbL873MNlI587b1/AzTG4uzops2QyoI4Ncz8yaTL
4lHvcI2Hk1u+XfsMtOO8tVifga0bInYONeZeUfslY95pyPSb7sCkbRqn/73PvjwT
C8OqZwCHpbxgEOkzm/MKhTOk1cVQo6hU1eHxyaDG8oU8NzoBiXy9zFw0wmUIBfm4
ibz8AT5RuYPToU2j3ZTG5wAouO2OWKwPgjC+o3PGhHKDf0gxWmgtvLsDVTxTAXND
IMzEpab+py2CR42MPh8tv/gDFk+Z+82hWNiT0SlRiYqUhEXiPY+YGvnoHJQBG85I
5oIeBbBINYYVr3pZapdvhju9UcHNTSxiSUo/QPhKIsa0pAvdAQAV6ZZe6+wMXV0Y
YxfKjwSdYIOD8Ei1x1j+SHFJ+WZWpZBfUygkWTP55nq5NpnfJDKxkHQiaS8UyjvB
YfcQekSk4JjiFMd07mBP6zhQ8WusZD1SwJKw3SNC7BTuUDWQXjp8B9vKUXQKjHP+
O/O1ww6at+DPYd6ME3YcWU7xdSqSHQSfTmaHt5R9Fv2WAxc7jDcLVDgoXGVg3txL
NbDrawB73SZdgGjzuZ/DQKOmJt5OQoRbIHXT3ff9xk3EuwJxyEESsD/nwN5WZkul
lM8cdaV/Ii/E41nubkw2cCIQN+X8DmE22vWI3XOLuNkhhd9mGEgEOKpYd+fO43ek
9eTU9NI9c09BER+d9JEX1IPOeynNEPH3+2N2dSzgTaYkuqkQDDgSRR5PaR9duS9J
B+qm1hN4Y7OpIUTKb7yl6hpV3bj931gLmqeUIHOexBrNG5onZv+t6KoJJTpbyhVj
SxKZrHJQgEcrkxd9GVQa8CeLc1o455n6dFErjKfNjeMiQa5AnVCAOvV4aH6CNmo9
hl7eM94QW9nL5D+7ZT8iwXdMMEYSBoLyxzCN5aItez4qzNnN5QjOAFPYkgisURMG
GdV/kPFz9WEp11K0FFv6kdYfXkzoyQTR2WFflyre7O/nrrgit2eBhva5KbK++f8j
+KeC/a2iSk1ibMbt3hlKegTeIAB+WUmY/GUjrn7LoW266Tkr4uKzYqX8slaAd1jp
3eG4ADMcEGjRJWcEuE70y5TuLBEtTy0/xFvE5BjMcZ2hX/8FBopIeS8kzHBysg/X
FXkFfvM+l+yDVTaLcKnxF8YNoFy7JC+moPetjIHaLYzFxRULnK6GbbmtNlfwwJKH
nYC8p9CJpS1cm06n00WH98DFWm4lvaefp/WmEPAwC3c+pcN4O/FjPqGnA9EWhOGB
aiMI1O0NmPMVgfY6/uP8LfBDe9S5b3V4NlB0qle27g/eoQBb5iM0SIDqhShYu+A8
O3M2APSmwBethAR0ow4lCCP1Rd9X9j+CHLc1IIN9zuOEtSTnouif/0SIAQZdasWQ
udbUmrHpV+jeZD9Nzk2ClZ65al5U07v9+r5UNv/TH13jrqAhLyOpj5hEYpgF57Kf
tRfRZC11PoLpk8Z3zmcp4HiOdipIzvsxVhbHDrMhSB7iCfYIJX0gsrBMJmOH8M31
K+y+DJI28X+psxgExN5LEOxGv3OhWzd38QTkdLGPVcU2eDLrHo/Oo58BAaWmXFJR
g5vHcoNBztXlPVm1auwJXiNYLPNPBy8okosPSSu64BC96N2Y/XKoSZESP1Jsko3b
kh8mkc6R0Ku+IwkkXYgeysZBA96w7GBvddy/0p643OQJ/n8gL2MgNKHtEdXd3fsF
D8/tfLQ03MkXwYG3JHpoLlpN6YPXaft+HszsGkWHHSAVu2Qxddy9lPBP2wJa7sCk
Sw9n09G7oKTiFPTIX9oFqJ4lfEVOgFWQBKOK6J/pD9m4JirZoEtA1vJbmku33u+3
R4i6A9wtmjNF3J8MdoKmrMPt07k2jAS/Tirea2IB4nH0VtTSmSwN0FpI87bKbHhG
tj/KeJBB63SrjA+IIO8sV3rRm/+BpjuFxNy8u8l0Xc1qQrXTAgNZAGzmQEabCXcj
v3xOfRIN3RIQVOPW0YFTMq3eBMlzWCMrUkedtP/Q18CMzU1XtPc8T1n1fDpaG2zc
hh1iscr4p7XLCfTAX+ezV9iN8yOmcGfoXMz8cD0nSqCpTCgtS2/VvrZaPtVJnbKz
3WBc7csXfXfz0FhiT2SkOY6wcL1DKY+aj84bpzdcZ0iQSQ0OWO3n+66cFe87FlwJ
nL+BZLBVSc2fhNjlrhtcGDTZp0gxgDLiQWs/a9e5n9lIEioWiSGIeSaVFYp2x3LN
DTz3FRB7/xihcGD9kh+2bMYX5nrAQz3JRhOD6Aa3Etp0LpwilHGzP8NJFinE4Lsr
1V8sKoyfWbvOdnzjB5jjybK46vG50o0FpMI7zCDFpuAylpW1ZyQe+hnytdggbGXb
olrpBvGnT8ZrviG/SEqPMWU7FaO2ABC+i/CWrLShyrMWK6OKiQ0BFfe50qMRay+v
dNi0GtDyKTQQawlEG2jU3w395xz9q9vB5DNB03o9iGbo3yoL/WZBUqyecvF3ioYW
KblXKw51gkgFBR1rrcIN8Ary8qERbYhNxW0SG4+g9bi/DNKaV1QMmpIEhCy+J7qO
Qm+k/1oSUVRQTQfLqA2Yffkc1ayV7txzUpe8ygC5o5L81eu7qX5C4BZxSbtcpJPb
RtFMRWGzN+E4DPFkDZc+d6uEK7qaktQmfTjliehlerIOdSQA7dLWJHY+LfT8MaUK
A0r9vpxIk6/dWmRH4G3eEd3dxxMXEiknj8+Thg0Fb9ZEVF5IpgvVV53d/AAHL2sH
QZ4Y1tqqJnLUheEXtgkiOR8XD40GX6kn0MeWHdp5kmctsjmhaTIiyfKxEHzSL0st
+Hlr0BY3I1qF+QhU8DiXSUkIOzpqxuds4/AMTdFdL1l+nEyy+8MaKXpPApl/WTjz
bZRBtl14yzNgBKLo08/l/WAOAbRoGs3voL39DZiHuO/J+jNGvhsbjLOVPPwWGHYA
K7p4CT/hYT7vXnt5ePZXTII3/hEFKZ9oJawHWyjHL0fzgu2r48Wx1YM0MimUO9BL
+T925L9U8g1duM/L0GqdW6HDL6JcAiJ+OefMVUL7AaKdLZG/Rr3NKFOD08wNaz/u
dST0SNyQS5pIoUNUNCpdjbcV5uwAnHI5KraSD3T8Z2sdQSVgox+enLdt9PCVIIe4
v3O6YozbN5eK3CE1XIEKCl+jvWboVerwGyFgvHWDaHDtUxaRWFPYppdCgAnI2LyL
BqBrb/i/2a/tWjv/HzmvZar6r8StvYx0a9zNFS2a9PdcdmkIPS4TLpVy00JxvJi0
RXrgBNflwBVtpTKHl69/JMfe8xph9ysV4CgpMEQERJp8sP1fmrxDqDgcxelSHc6d
reWmMJr4znk4PpietTfdWr52Eiw+VaJsXnD0xbbgpcJOg4vjsMKN76PsOxzebct/
dZf6EQLvH94DZTkmw4sb9cz/KDpIaJDslB+QezZoJ2w/IKd/Jzz97msxlizlJzHk
H+ATXqZC57Es3VVkRh/QgftRBPdAaa3UQ6cad7nmAGUUFptMujMofyOnBMEoPNzW
Ngd4Pq5wr23baCZcnkT4+voaCTevjN2aDIaDOy+mPtiSi6oqZawLl1q/XPI2bBFG
9evnl1PmptlJCJ1LSyy5NOnOkV4STNxNs8LctDwEtSgGHg6uceVj+fr2L9KKHS85
lNZdlT1zZuBCaQVmi95Qk7topf0ANc3uDW+qeOWekgU13ez9k8kHb+8vRAQSIPy3
6L89qpx2TPPi0N4e2SMurkLq61I7R5W2j4OLNBcVyqGzPuA1Tz/VjgWRYFTEiMRO
1UJurY97KaarTKAyRv/eLaZ0d/mUDGNV6PbfjvV0amtI1gPqFLE1HiHG4LEVMNFy
wbfKuJM6oRSXy8W9xQG48v340BR2KBx0T0XUetPhzFLi2alLiY4peoSyVSoC57AP
/t1+8Nm5vya7TbA2TsDiQgc18FvxbWMll9xzKf/RuBhpdE9oUXI8xSR8+3Uzq8Xg
AOrMfJa1nct8agZ8MY2WlLrmBbFXDgyx7719Q9LhWEHtwa4ZinU2hcOu7kbA+VuJ
VJRhQGNilZyHLzC3EAF/pi5ZhfsJaFwhagzKUG/3FumPWtS+XpX5xfa/rFCN7BbD
bvyOVj6PEEcBE4O67o62TimPewDyfWDodzTKkakWl9uXgiqGvMH3aRrMMqyfRJVx
S+I9iOGDGsXWPClUNLaQlMG0HrArx2hxYsshWWJk3ZNuxQdOU5bmNADRLxDk/PoQ
LLf/WNenSK58mdTb3L1ycXtkLYa/lU0lgXMA872mwqX98iUnmI1YFiNv76cOmpni
+jN2beUWJJjkBowpDZBC52dq0/nAwdVIznULB2U24BT8Iih5s7cQhhCdJeauTE+U
OKgpynclPN9M0JoFSje4oY3buJ2M9qPB13sXItk2kPxRWTAf3Q0x240DqjyNtaV0
KXvq5eCyC9EbD7y1aimi/P0FWd93pLv5LnXFboaWMYDFP4LGMadjShFeB13N9apu
EdqBIzDenF/uLaQYyPS0wAB4EWjOhXVGuOaLazy8rdGblzINMIxW2ozkpR2urlzX
Bfq+ow4Z2Kvo8Yqz1+PB2mPqaASeMWz/zbcwzYyx2SVg5D/mRaQy0KwmRUPW7FiJ
q+s4IvQjJ+T0VvkyaPqRAlYGHkwvLoO7mZn8MJDVjdLJrwnnX9oilHuUdjWymXQu
3Q3WCbvH/aoB0W6+NNIeqnB2FqPQ5tHYC4+4WLmY4AO34VIYXSs4dILxfJTEo7ra
ycaXC9ic3QNVjmWnLyQAHGwRuX3bytJ1IsCHjcTlU2Uyxm3c4P7nhBgem/wNaSjk
wxlzSZHATEfcvn0nPmT7Z98fHBPAgmYE97d/B22wZBCCrfYwhqk1bCDEUl1tYXvF
4nGLrPg2wkGVWJ9Lt44r5dlC9nzdoWCx34sXbhbacAl/pg+j9Zld+RcHnC0JFLR8
be7hilgRujZqXflFou42cIsV91K2Ns+LdCnTAQS/IoHrGd0yj/6L4ucd3AwvdSYy
/bO28fG+cnoBjnvr+lf6LQOjDzdro1WE9eHoGGR7bFikM2Vmueh5nzcTWROriWpA
2XBPbAYcBE9SETSeFDV9+A6dlfkuMfVsmOPTiUXE04HX6G7FRth8lpMkp5yG8avG
hcWGyM2pJ3iPqyGmA9hFxlrQn2ZHB8PNAZWO0vVUPPGANd1G96D5RGeoeFmnfwwT
GV+uB+f+GPKSrmEqFgCTuz3LCl1iRuRODoJZEJ6KIO5rbdLJ7B9hRu7YCsq0dLHk
vUEr/PxyL7a+hwHE52ylUqMK0k06jIEH2UCydoN+zzdfkXrM1qwbWXltxACvdLyy
kHiHcJpuigE5+hqjNPa1swG/xiM9tzbL12k3vFe3OwIDMiTiQ3tq8myZldnCHDhI
XcZrEBGlOSEpqvbf55xfVHbeb68jyRndzAFzQrsldCKoG01qVERrpbcJJiQ0AJQl
TgWGewREs2k+KxsZlAO51brq/158c2ae3M3e6qKDT0O41A9eCZcRzRTvyPybXVnC
htud/tznlCsLJbDLrn8hqo8qVxkc1YjIEAvnJ30oTpt+VAQUfVErxOuViynrQhGe
WRSULJKfi5oeKvvKBdxsRFp4GxCx3UQzsL7AcntZAaOuZJsY+OqC/VdrY4kNil04
feLcFDUDANGWx74BY4f1XO358QgNOng/tdy4pQKqzULagQ/2KVKZ22Sl/TeyetFK
H7MGjTfKWeCknV8IZXbVQ52OT3qVN/AwY48JxcsSMcIGYuV9m4trPkH4gthCWp95
ogIhA4YjG3v/RcPMsyJs6J/57Qk4K9fGdnmR4KxSSnN5/Lx7KpOf3APPnfs1ljF3
HZ3Hpi2qsLWnlGtFzYjzg6GdDTrKTars8ZDTERQdtQN7YkQqX488JFfhPqv37pmG
EnPh1RVD30EOkmut4nVaC9WFK2GvUxRHpUb4zgGNEnw7quxAje+AhROux27zjWwK
o38K0vrVLiDDOFzJwMM+5Udq/u4SpeB68I3lzD8n5IVhdrjOOFRd29O5ECRMxIqT
HEquNnNmmpk/dR6DVb6u4tgGte1ZUtZVutgBInkdHa3v7/q5OhEBj6SsPPRnUlcK
OfOLBdPjeCsrRsnYWS+5DFjihbV/SocZEKvpI/YPe6cckpBBcYP3hIfh+imbdjPe
NxZudJDw/WgIRa2iaFQuv3dh1mWQMc/oG8MRIJOGeFBRF6+c2FQgL5LGIHaSoxxh
3wKYlp4vn9yV0lgeHq8AojkbkQkw4iWsdiTWlhW/3Sn3ZYoCJnfDnltMEgHJYbeb
/o6ollpGL54plBS8mv2g9kwUMnodZ/6oxtLI/LDpmRHOkWqbvDjfvZkWiG1O8k/b
aGWwBHq3Affcfk/oV2XBOpFHxTCCk8t8s/19D7OoDz/Dx+DgfuDyEK3NfP+XfMrM
pde1O9Ew9zGNoDHMFhYNm/yppX0H7G3W/VhXheYgGp8WVw85pmZsJGDkCLwfg7cc
p3TTQGQhvoRezdI2xLTKQOgr4i1FDlY+8heXwMMzMZU08f9xB++aNtpOk+8voTI0
HmTg0yBAEXU6AYGzDqO2VkkObGd2U6QSuVx5NFC4XePG6mXjb3kCh3mimZ1VDXc4
5h6ZGOUYmTQpvUkDzY+ZALhFuYtQjVLyLtKpAbzTu4PNM2gim7xjTUUdMmcbMYfm
g322a3tmoRb561iXgZFJW4csQck74IFzkN9h2T98PNBmGFbLG9oZYTMb3MpQnDmG
8qrz1NGoZYtxWRk7QuqrQEQMERxOs3H57kr0YlIc0fv6knmkK7ixlbKAcw/X0yXf
yJAxavGqr7arberHUDZXnDL0G107Hw81eyigT/ojxE2LhVC+zNSqpzvslIMmBawE
MnniClTB58dMDjWpuNC3u81HuCWrJ3h46MfrdFUUAXD3GiaHtTT3OopsZUBubY/f
0xY7SGoj/cMEkMV/xaL/aXgrpTWQcDbAWxzpzUPFfPKq6KAKjSFlZf79WP+TvMhP
CdMb9jM434sD1Tz9MpIvPGsqwwzO5NV1Z1+d/Td0euY0m+ONKPI3kHbad1N94dog
zJ3rsb7P8e15Gicvch+xYfSObAd2+YbcYbF5KpoTlURPpKJD8FHGZbC9uFsyLTH/
i0ChFMQJ6D/aNG/Y//TLYZejr8hWo+O0sBu4dWNAQxEV3q7eIr/TxE+yOFRiDteV
wRSQLwkPTTzB6eS9QBstmKAbi6A6JG546J3VWfPBEHeLEKtuNC5wU/wcy1b7NqYS
YxNYQ6fsW1kmz4BxhIDOUUNfaAADYTfwPn58733dDGClLmACMjR4HyMirNCKcGxn
CtjV9C+ZrEoqMlo2qIDcsA1BuRQ+5flZOsuiCJaEkie0bCyQFRHwneeJcxvdW9bc
WMcGZBpSXY8OpDlwppseIZefH9rP3IZe9fxHqSDet7FmHYs10007XkDB6wyFzHjB
HyC70hPY0BsYYEqa4WJtjEibuhRLxImNkx2NCdygFxkX2ANNqtEbVSFQSZekWR9y
zEYkzSmkslIN3VhMsyYzUjkgqmRPGEcKyG/XZA0YxibFbfl7ZBIZc1J6nzvnLHZo
VfHatpwH46fpMUqWiL3Fr37N3lnwn97ZwDs9Jwg2CMuM+PGCiEj5Xz8FIsb6PD37
DAf66lSeWxWzQToZ2qyG7zQc69/u2JCsRmZOTgFAh2iHxFAhhzrz6WFl9eEzaIje
LVQrdkUBBQYNTYjchia+SHyEJZ/N/DBHAWDHkIsg2ydsTOqOUvODU4A802K10YD8
wdF/euJXa5FFCsZZLsOp5rzTqbCNTYBbP2KrxXfFNA9T2isHMU3Kr5ELghGQhTZ1
6J/Iv5a4Jy+0XLaiIeZcXrSxNv7+D00fZRgFScGXFwj7ysdQ06pkfFgjw5HwgRob
8TV4m3pUlf07Zbr70IWgbKLVdF4o4VDnaQ+Xpy2XF52PC8ynRS1JCYW8aw3YsYTS
r6L7eeRXjlPGSudwHoEi68SRFY5PkXlri0iqEmfhOEDKFMViKEQfRxbl+HLNT3Y4
P6oj3yKsT7FeTfUpSwUbRKKgY1xfAtFo+vdwX74scCwJCeSp0VFfXZkqX/mSbUEO
VvcgM1KlnzM5F0SdF/AXMQcvhtd3N/HCQe4T9j1u0a1she/BFf69MFsGvze1XftU
Aj4ygaC64FxAOpVwCZ4Id48CX1WhzRNby9THxCcSocEXOcpwvtCDTWkp5P0NrAEe
rB6qdFjQKbhv9VHYNXhe15LB4B75Fift53m2rZqYm0+6h61B9QV6sAvT5ks7HWMX
vcHTEIhwqzOgjK7dlCkdF/cDrrBmfHRlVCvLfLsBZlxyp3CkEs7i9KGyxL9QbpNl
u/Or9u56nxgHreoMSatmwTA8R7bUn0Yu5kf9w6+ZRRLNkjnkFuKaNVadNuy6oM4c
qjYrPxq/5U8MFfoniGYr23JBgcmQmJ4W+qtiETCIUoq4nlZ6iWbSRA0JQ7puHjK7
M6ZIvU7wXim2eQe4l9+g2ShDJ8HnyKGLFgbZlZVl3St8PeC6wv60q3unfIddkmT6
5VeEt2jo0j1vZDoqZd4K0yOH1P5j01kM3sG2mjh2GDyF+5Tte05uAvu8CgxEy1TG
0+R3p2ND6kC3/nZppK5MisGieDH8NyOaMOD75/gimgb6P0T28svqgcAnQfmuVMX0
+otpAmFTR69FxFo1l7FjAt4S7xuDyO0BydIij8LB6+iwPgEz27moxVA4JYyhUk4s
VBj9l6DEpzaI+2EmUERJgpyToMFcaNhSnTKx7FU6wfyJUUq/Fl9Foa4F+cKCMnXZ
ehGTJKXoKNLC4FkHBfY3zMqB57uycNgL/eD/d35vAK5pVWLq2vRuWg/GlUEvVlkM
xvv/16autkvdFOZBogbSCMzNotD02vGABnyc/0ldMLnOuU0GxJCO40wDf+i/T5s3
qUlQsbOxM8z+qA4GK85ZreeAlz0f4aOWo1NwA5wIbnWPMSB4pC2iChYhMCf20emG
cr/IJt9AN0vj5TU5laFIggQUJ5UbkiEQwaTQxeDglskCfOIX+9+E6BorhDUVlpGU
CRFQRjitP/50ZNrr9q1RxycHU4YuxOJ7g3NosqfxpOVU173A00aHgC9TP50EA+dR
uPnytLcINaPUmpYR4eippmgssZR7fbdrCIIHUN5WFFbxA94XTjVfvpVz3UYTndBC
crRH5jj2R96vQrPnhOSLRZ/pxxk02VhtuLxhcKg5Q4khA/i6UanmL8cwAIibzQKF
Rs3Vq+vodSgJ+yKGTSd8JT6LMfpF0qNZ7Wl+DsHo/5F1GKT+Zqg0ey4I6/AGDaBA
6SPauhmKbhqBldz8wohrVesf2yMJ+P5d26aTm5Zd3lD0EaDM1WAiv7GmgnjuBVDB
f16EiULNz/uCEZP7I+RaZgU3V/73XH8uv6JdagoSuGi3dFeTsyJkBXbAr3VOBksy
QcTdL9JOLIuK5GL3Dh8XLYNBUso6DkWWq8IyXyKOAmSuwtAqTFAAJEoAftddMkWI
GuZQRrepfNDRC+89Cpl9epFO5aQdWoxrinZlDSI4ErsEESqZ9BcW9BSTnPc1er6s
NwqE58+s5kUDDDVQou+fDD79WgXH2kgNc5Zqei9kfvsebojV3KST8+tRiBI+D8z6
+eHOavKsCRhi8gCOQWj+sqXtg7bai4SBhTKXDwFPhIGpwshOez0tNVtTKaomsYdc
xZYuzHJ0nNJyaYikQJM1MT9zoIu6R4xtyoj7EwpUbvr+iBC04EkJBSqwf7LK9sgk
7i7/elO5C5zyksiAGqongR1yI7VUHqMIjZwpdAibstVJhxrW5XJOQhbhIgmnQk06
tddrAsrLo3IcuzcXAeRpU82jjRJkqNb8ZWZBnbKWa8kT8z8yxj+sjtEQcBWwIiVW
iIVETIQW2XikjbMHQcla4I49NfzxqcDo8D30uvfPdvbzrB3Q5OuTbEcENN65fbib
pec+KexXbybzopbLOvQ7hmdEwF++HINyO2WWP77l16PHt9HNSmu4mgEsOp738CGU
wPWcxaXvTGXVldqNfFHqrYU1VZNoJIaaSALK/KLs4GF+XKBdkgM5cIL41ud44wtf
A3ljKehYL80YNJpGMv5XbZFDiH8ULiwiLAAG6PT+w3AePcqHf8Dc5AMHjzbiekyR
GZ2lGZVOQhBXZcSSggPe/Qf3QIao7ccac+Iu266jp1GG2aD2jqKWm7AOg5OlEC3Z
qzPP/3RAB3Z4G8AYFNNHIM0QdR7BO+Bxp6w7PTOAo2Z2O8yGZskj0LRiomSQRCt9
dk9t0RSdBnRhPl4Pcf3QRkqPHJee7YGf/Nr+8RUNpBSl1X4XpYHMmaFs6lrW4isF
6iK67HoOy/kRmBGh6+yOZuPrvBWmoF0QzUZnXnqITX4VtY1RnD7ZhCZA8JffjqWn
f2VbY4ivIWd44k7LQONxPEeRGp6SIFu8/BqU5OWQct/xnPkTlV0/G3YW8+YMgNmK
HvyHNswMRU43we1iW4x07u3SBAr4ZSf6n2lEjuuBi0Yy7kErBcm1k945FkH4TFlf
Md/r/bdOKLLtcepBPmfMTnNCH9DLMdVowOgYTHi/gORIdH+nIof0YQz5SjRb/KCX
LSobCzKil52hPk8My9S4FyrfEYXtssj6bEk9AFhdQgCawPDDa87og2KoD5I1qYiG
kQKiI0dPfYGbWC65jJ8GhOuCZ0Ee8nA1YhJ7ZOMpbzKTVT5gBZ7sztcZHec/pIyl
gU8Qx6PrhCi40chsyrI2wB0Kw2cGaYOgZWnVS8bJAFuJG3H/iNEk/kWgW6UWXkfc
elGiGtA+Kz3IQXhu5nsLJA1CGTb1zWsE3WpYrFyxUwJFzjBVDGl2d+JV2XoEjN8i
OXb+JFRqxbedEHq2YRyOBnn2tlRgy1U21/y0MjQe3ch4doE0i1RoOkRa+l3OoaHB
3U57By/cTP/fY276wABKNpKieq67hUUMfSitCmWME1QZ+c+kuuWLzburaPSV+oEr
D7efixUAUwS02SM/abooQpmB+b9bxygffie0Yhkpddz4RxkshS3fki7dCNJx4Yl6
zJ8baFqNyaRkSPoFWfnwAsnIFbmzgJgjGBie4+UcW76327mmf1U0TmIsJL9P8/wD
ZgUpNRs/MR2gbMVrFhKspI02UOWM20xxSz5RcWYp7XmzlJSlTiCH+qn2ulr4B52p
hpgIKJVhhyNnO8IUi98mfbUosP9RMcCI4IQrfCkgdqu3BZTkoOWeUss12yuu2k0D
9dN+c4V2X/MKCjEOh9ToBKTBDxfv3eWCkHD69yTW1EWJOjJM3Gr0MxWZdduRgbV+
iGCj9LRJ7uOi/s4bPR+NxBnOK0Y5K8FNttlPzK1KghYDr1dhl9p4slGRtgQe0cks
L2iY0NSYgnqFJ40PUtWTHWBCwJgV8Pc7MChlbKJGOCtq05VFx5P6/bhdnwbmrpB3
RkhaH0jrArY4tLasZZAbfA1pnJBxCzwefcbUysrLbhyWI+piVokUTCuDPconL1nJ
CJUtfyyz/KJtSKLe5s2sR/LSwDVK5EDMJJIQAwHFHCJrYix+0UHDgwiz4r7L9jT0
/diV4aWgZEBjWf/OaNqlPyqP/MtjlWapGq63DkvIPTKBn5Xsu7cqEk2Z6GtI5NCd
w6oTV/6XRvz2FHoUoebNnoXM/O1t1LdXE+Dz1ohgsPxthnuPqYHLem9Ghsd93vLj
NFZBVPyPF91c/fd4u2W8NzWgZGvs8ZkUwj/26jkRJzV2quPxHwKc7ihJARfHCy+m
5NDsNq5Woy9lgf0XJKk8cJNhA4l63Tv7qruEU+iF07JQeGj3YTlAy0Cirg7vkngG
PKU/Mx71lluJvXBkSmS24KHLspJdnMUdXnizZdy27/KXaxSqEbQWeoBranD1i56B
V95zoNTHqna9tCuxA1pQQBT8566pYUAaQRXMXMz71gOeMvUHoobgB4Fko3pAhD8H
pKY4rNemW2CLQQEHMjUCs8zRyxZE7At0e7EJCAZW/c1JVh4/Mv/P+P1oqDObBuNR
7pK1YAQxQe9hbprxISr4UMo4jVN4EzsWInaDVmvTu3GSjWE4S3/SWlmDBYuFSq75
nppDJrJyI9mu+N/QmoxSo6HTRuwQYaOoAwjQxdhy4M+qeFexFG69uvIkVewKfLH0
gph/0y8d0ZXVXMhx84SBESVS/Q0c6tEk3mQ4grivw8FLX5fi6jZwpG28GVk4Us/9
GY71v6a6kwhRUs0y8kaThtTKy79zS5NmWVJS6cwtva2hdaHdRyhsqdPppNdoC9QR
MEbYddmBLHk52yZOfmDbOGgZuthee4RQhBZG8fb7pY3hbXRZjomC6glfJ7ENiz64
nnnHhOkWYKtAx8UD2sxTzy+yWvrFxlYENkF5nEHjhwXLXDyhBej7tr3TiTGx+qlj
B6yySrPVb9KKvqMy6nX/IOCYKVcImDOBgBXcov+LSzs/ErYk8XXyj5jTcSDRE9Gj
g2YFYJTTuf+0HTI+Sb74Y3vwYYxIc6RPHUmtimD8+I6YPx2JudpON19BLuotBEJj
8HWG4rQmwb7ezFVLmEN7lvLfoRD2okt+fDaynB3bGZVLYMScpkVg01VW9TUdWujB
AgESCho5Tm0CUrM+n+/B7OneJXiyIXe8Zpvo59+cphHfoE4gAKfOMpTUkUcxtrcN
n8Gz5oLrGxSEQ5Qt403GBu8NKY4Ql1tBvBYchdlA0MGU7h60Okfwq6PLn8ZwDHaF
2guP/tAIcgslsTSECODkEeGZ+FL8TlR4ag6Mj5FQ69zyEbDlT8+dPMXwClyAVh4I
lSkv6jlREYFUkHquacbwQWWUckrDoYD3kbz7Xv0xptEU72ejiwmLGuF2eF8YlZ7w
R8KbgQNrRWbNV7l9QBch6YzlME0f5KYDSfoEU5/9bpRQM2Vl2hjNIOr8YA5qO0F/
xE1DkHMcMY0aHyMS7i3rO5S+e+fIHp64KyeB+FA5Q48a1vPcVcL4dfZ0vGBSdkC5
0sai2/RCb2qYOge07WUbXSnz8oh3lkvzAs0iE5IqChJblTv+CcKC1GmbwOWXpNS1
6N2xqYdLmsguw92xBYU2Tso/dMW+EMS4y6MsvQR4qf4v4tig/4U/pxYgf0J4O4eF
za47PVk2r16rNpELeSYQya+Vpa+6qgwLffIq+jm7fOoxavw8E8d3shb6Ob1Wzmot
ULpmpjNJQKPCduZ/g0pSA0z/f47Z30Nwg1pogP1a3FkEbPiPuXaJqHcAxCsOgR7X
WnmEEb2BUHBZ2qxCaXkD5z+4X+/O0p8mRmsxorgBAtMKbX+YanqsJAQ98DU3xWlv
X4/kvt7XiO4yVMV3iZSffZwe5OR4hOERVjJI7yxqaRxlZcfExAZHz2eC/J7Mc7WW
gZ4LtNAanB4dQTzshGsPvPrHIZCSnQF3Jzk36HdeEhfjpHvK641os1QzIH9U459j
tNZKpPJvplUVAKBk99weTEf4C78ptQ+nCcPlqc4RF0/AvNmmXhgdtUgyuSyiE1SA
fIqViDF/+dtUpmGizytpmjuTxN08AMsYusmgS07D2GjoAX33Hj5xsHMzNKW0ugTz
oRHkU4b+0EEwnWvlPb2GAkWZys0jXd0zn3DDCyiHnqsjtgmlS8/A+gIEwxWvLgLZ
cQX60PkYvDLL7BqpUSJ7NlPgGGVly4YMeKmM832e7qhb5ES/HLlJkc3CDxh5SheY
/v5H2Sp3D7EXLWsNH8uj2mtA9vZRizpLQptQ1xyvaNFX7/nyjDpm6Yee63VExqO8
Ohc4pj7GEBRBfF9nRMcH00mFdthSfdMOOJh91Ow6pAhmbdi9zl3CyR15wZRqXkWm
ubxro5Kem135SHAe43C/raoomEKCkMvbcRgD63p98gxDeOcY340Qn/DLWcBh6nEX
X8NCkKkmqG+7fd6hP3aewOnEMhEaoeWWSWcWRmhJsvH2qbJHvtz1JRCCjESzcj0G
l9pkY8WsiY3Z+VREVpUGcrRypF6kW3OHPYjV6xNkmQ4=
`protect END_PROTECTED
