`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9dIsJp6TbyfnEXvBz1Cko63jC71bW72jf9M/vtu8K1+8my8q74vnHGlPSOxdjXC1
NkoKUdUXISjXwCTRgfusuW9eZK+wYf267gN2hJ1c5G6iAyOwks7lHQj7bDUdKgAA
7usMkZhzuZxsBwjaMpE9v/VbQ6feCaN1WJvxuHCjEFBWMg+MPTXz4U1FmMn3NH4F
btzGMyiR2fxRoElBxOFrRf0RB8MCHfzbXr5J+M8VFKvHy2pkpZasNngNv4OM0yTM
eFW7Ohf7Hc43Z9oYi1XjuKWBHx7210wVB2Dp1Mn8fgR+avso5MD1Kkkk3yWnr6I9
dj1BPpdRhyPklPhDu1XkWp9LczW9nYEM46wfIWhjm5DuQsn+px69DeP6SVZLx43g
c3kBMwgPiyV6HCz8HBOOBGPPCXJhzMI/e7xBmR+TM8Hz02kIClkrmf1xGAxRifzT
SgjcQBEpuSt5Gvdt34yx4n1CzeAMWISX8caEzVMJvr4=
`protect END_PROTECTED
