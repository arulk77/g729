`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MsWppQwSU6wlVIR11FdZ9wagH2mrZdTqtB8BuIsuOurzoCUEZ5VE8Hyj03JdS+ru
Hx7fJV2+fq3G9JemFMwI9Ow676SS4BJAEuKdj3qmDpHVNCN/e++LkXzqiyffed+y
QRGDaPna75W5XQuRjaryX+nb7R4syU3oQ7q+VIzI+tH/I5JxjcEVtY1vrqnRVaj4
B1QW2IjlREYAlqUencIeVfUfhd0ks/m/NSJnreXxumE8q/5GKuHcvigNBhWd5z3E
uMKImTtwfcAqL20y6BDeYDzZektdtUfJTKu+iqvKluYCL5nFdlpZebk9GJSUFxCy
Yxah7+WkxTOXGrHEI62n2KU/noU9X1d1W7P3wl1NZ7gnyeixbRqvsRVzXA1aCn7D
YXIqXWokdT3g0rSMuv8y+wDKMWPRomltoGsb/FoD3blaJ43+fQ+4VfH2/fsxTwQL
25T6xEWg7bj5JkIYK6q+yYKUn/tNl1X0qsfiQFHM/7b26kqx0GSzcSkXNCI4s2Pv
7GjIpIQ4h17alOMeiTpIlA/zB5iGoFoFKU7Mx4HfFqv8uN6wHV450TH8RUB5uu7+
kXI35vbk6K5XrGmkyOg5gkRpaNxXsVUoUwYGcfPZjrxRxNeHuJEvRPx42SPN2lJn
iZbHfWne94b4qxxvEm4I1DiAyvV73e14eBu7oIxYxvG76B89ivAXcNrGA/8+uWnx
BKreQ69vdQzd6VbyDFQINw+FYdJxXdGvnq/NTGUQzJ5PXbjXDherYVe22RT/+tJh
1DSZFWCldTA4wrIvPvZ0bGUwO1iNW2ASRPyqT7uXawP26BilK8C/6maTa90OpGFR
MaUb9q1/51qQ28wgkZoMvERsBFrGx4LnpEyQssMjn2bHJE3e3HwR0mCeAFra2eka
wtInuy8uU4gAEtLCU1trOCpBXmBJn26kkq+kvdmUDJYyfYCs6o+tz2hMNZVyOcZ/
P8rr47O5Nu174NqFyASAfKRRXMpJHY+NnIiIxbhKgNZeANUXr3NB7+rDz/kDRHRo
nYal8PePNJEgFeGSUtwS+sxlzrlsFpEqwxVN8X5OdrcPwGqiy6UdbiVCdRzNmfo6
uE5xASWvkUlgmtkwMhr/AnU0v1sTJfqY8Y5h2eSnrl6DvHBy5Pm1k1z+Z2c7wSS+
b5VeQVJOiDzxcVYQH93EBQuOZbyUVEUbSfp0oRPhZz6SV8+xtFWTVCZChVT9xBPu
FyA+yPB2A+PWRegwBh1Vr4rBCt5FixpOaZ8yVNtlfQg=
`protect END_PROTECTED
