`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF45lm+KEIUd2Og/zgjn6duD/8Y2JhqIktBCrdj/YqlE
68UfV0g+CR3+DtsrC8xw765wHep3dV+hA/Ldll6hXcIrFwK1X+bab06C8nQ/frHk
dFsgKQQo/42Rkzty8YOlRDUUyZ3UeyPeH/Ccbh89QxIJpEq2ctCJ0RRNgVpa4bDP
8cBrrEKvel8W4w4RPnmOM+CrFQvqlJnfPpXHl4w4ilow+EPc96+j1kF2X0SFirtI
`protect END_PROTECTED
