`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCXJyIVwQ8DjqMlu5sOW5g2GagA+ialm7cEBSY2tP1aX
w4gEuVjA4bYdWVj2t7et+x+JMCxBpO9v/+xif+s8RFZ+k1PNciMVjGb53pKoa0Mg
qqvb+LRKaeOYejYOO6toWO9ryuKLg0lQk3PnvAeRCzt/7J2nZN82IIDGomr4jKfZ
30232zaXfxgtwgxYGzBvgsbJ8EyI18uH5SxJjZ08XFNM4he6OozaClhP4c8ge38o
RMOmtvHeBY4dwlAlgFFIeZSXnNvZHe7lwvLSWTQ8yQWTuiAaWLFGFKr/2buvchEM
y0SqSRfgQRZ1aQzwTmYQ/eDC6PwBkdXA8tCILoyghmR4vNy23XlUQHcInBVXFTBI
7c7Sw58JMwPN10KXoSsFcNY1UR2fE2+VjDNNWyELbK8cDqkSahLXJBMFeZRmMdRc
FTxLZBSzZDuHyxpqWbw09P8D5Dia7pJ+ojV/frNq9y+5CJMkV9j0Agn+jbVc/AAX
XhsgjryvINr5vBl3Iav3HRaF2tm2Lq6M8PqJrl9MYqOpwZEfG8Ak9lBCZKldSEve
ycC7sK3N/OKMtkvcYPM61PdbpHp90+q8GimFTMCGNoaYAf7mq99LtEQV2w4CxlWU
ftxeYl6t4iR0NPhJfqzwskyEl8STFyTJ8QWbCpgX8EIv2B8qQoDA7BnsHLuWQHng
eNRqvEV3sFHccF91gQW5VmuEjtT7f51hppzSGxXXGsq8kcdcoNmZOlntlkbrVnWl
NXTYQngF6aDu0KDisXUaCniN5HFTpbijDf/rOEVTMHj5fb9/KMXx0AJoaB2JlPk9
Gw/iWVnl+98kggbbk6G6K31cHgDe1FR7NJxI7iwNV/Y=
`protect END_PROTECTED
