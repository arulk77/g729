`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46bZHUqHnRAOwzINaesprF1P7qj+cVvayvfkFb/WGh/d
QzO1tW9XZsnSMbahhdi4OGVQCYwJkRLElTkijfsL7pM4plIQlAbAIZb+aVonZ1Ic
4eel0ch+pL4S1xze5qLu+i4D6Jaf0xy2kb+Hy+OsGOT7PhCRe1YHU909KWAePMub
Cn2DOOM/m9yk9tcy0aKu6+AXfIKUqdf+NHbNa3m55CA=
`protect END_PROTECTED
