`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48LvH7O2yf7rmO/vT3SsPqmj1BGl/Zv7L4KPVx4ox1t6
5kaQZKcoxUoKpBDccNUeVL1WltRwRugyqFzcGlsYhpmJVAkvr1weBzxAcKElaimf
WDtKMOageHfgk+B3/RtCrsv3DX7ByKy51ATdFaujSfTjO5rTFMY+QEk9Jo08R2a6
zexD27R+ToczZ9E8UpqwSbZxR6LVTxaSxfIh5ZQ7Pji6Ja1MegfOR7dMxegWEs6k
ubIm9utwXyuVsIcmwzfLxfyNc4e0TWU6L8bTunk99AP5WbsbSXK6uH9ZZleSGMvQ
f1+TZ6kP2ccwbCUD1AU6Wp6p08Coeyr8iYE2KPZgo9cCHKRDLwa+aQnHfUucLG6K
vagjn/I7zWVKDiG+1wARJg==
`protect END_PROTECTED
