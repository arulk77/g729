`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
yW+TrHqPVBe6aVyd16bfZO6pK+Op+JffCHta1wSI01+hvWfuwykBsDOfHqVO7EH6
8aSX3H7cp7Mj5xPYsw8pkVZAxwjDiNaooLtkgrqVF76nkbux6w26rCb0gN/rYdk7
+TPBy57YSabAxDsGrNhrmBp5D+V1biKon3RGgCQdg3iShLo8XkyWbs1WKTwMJ+8d
+1HN+D1oRSDrlqJgahCCu/iukR/HP/I/sagfemSH9lPVKe4jpcfpzbzgedXOFdNY
MUelN1uW74Q/adgSwhPBdlAJCWyNjYtOAOldmoKUGQO7SYXMukyUkTlkr2+Pl7Kw
Tkz8gNPzXOaBd1UnCdeMcRoAbQHOfcqYhjJKHPxRPEqCm2R8nTHcATkx6X7vkebj
GkLg0xZNBs03tabT5mzo44bjiOG1wykfrQHrDYDh+XFRykIpQ5lW62Uu4KXhlHFt
Rn8pAF1F+TBoiYOvnXyZ9qugeKhAYE15bYdrxAUuTeDuRLojQsFe8iwJUmzuMkv9
zuqzWPIxog9cG6yZwxkv6qlFt/qPW59Kv8pKf4MQQol1MLLax8b4owW3bHU5JvLK
6dDUXb15NDQrRarPEI+9b6rIGuErAhkvq0FfhON42BfJR0LlPVeVGYtHrYCKDERH
PWyw3GdMv480HbF2vmvk6g==
`protect END_PROTECTED
