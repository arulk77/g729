`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
u7LQP1vdIYwNq57HMHUx6lpLMjNLEFrjL+8iFImOEfUIeRFcbEet2a/rVvyTQxJ4
FMxvf7uJD6El1aektaLN0Oz0hiW9c9wR/BRtYqfjAu6D5+HzvCDwi3JMzEj6cZid
y1Prz2XkCIkul2D6qf0Nbdx5aN2MLkKf7lqwfZx+cFG6iOsutON+CAZCv3wZ09mw
mhLbBPgueiGorxJVUajr8mIJh8Wse7VHQ+bJ7NNLA1HkCuJnkcQbRhIXCjcBrrPC
/Qtn+Ko1cYpwDq/9gqk3CN0XAqz/v49moXYQn86XOJu55MWOPdvcqDfAd00lGXOJ
bHGvXFdeimYOjaT2+P31ZBW0lhRsvNLDN8GEbmQ767n7XapJZM2skskjDrWJtZTI
Imb33oRn57187VyQGvJs/QV9LxLyOGgkopIzJn5NokxfdVidHPtfOIhGBvOvwFj/
Wiy/t0X73ESRDxAweQMbAb2rJlUlzduLLtl/25X/bGKhhJhbNdN+vJUZYaz4+CA4
MKP1UlzRw2iVUYLTxD1TKhi78VnPl3g/N0BFY/D9kU1ZqXTb4rKU0o7pk/wTEXA8
4/Y8pS4irlM8c/bWAbPHGNut+vHxXyF+c74UzVdJNW3Yn1YHFZVZMAR1T62J1zmi
`protect END_PROTECTED
