`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMnBbaAKuQLtSF0w0s8qE+eDowtGYQCe5/KLE7oC64lZ
8xGBjZTkNrKL5snrzPRJQfc74X5TR5pHgFWgBm/IZ15CXK0L3lhzrGIubdU2LTf0
GNrhIqX+OJWIqdkClLoyOA1e9f2j3ihRf3HO77tmGKrK30E/Nrhub7Xx+aDI1jEU
MPaCr/xP9vxtRE/HbOtQ4LxXic+tfr6KhGWYBHDIOnCtsSLJn6SXlp6SXmge4tXQ
ezXhc/ZKub6A0lS63g+459brMi/lueF8oXMzLFHS8vOd14Mr9rDsPDusrjlTujjn
28usEFIVXNpeiLp8SQl8S6c+1AYkTNtfc2eWvC+ATLlvoV9V4F2Y2+MSiXlVT7Ir
TLIcPm2Y1gSdeOd5HrbcXoKXrhkh1A5Ri3X4iePea5dxHZlpAeyFdtcsmAnA+/GT
Z5jxm4UKES5lHGsekOSSU0pT6phmfFaPdeyOKOoycBEq1WiyR4vQmI4ZzXf8sL2R
3cL2ps0E2fg+wQYOWTZJtyIzIBybMgKIyXYNdonXwCLTgRHoTP2XGZMaTPKFGheJ
Y6D3/npklb5vfeuiTgTDpZ6SWfWmZBCruqF9zkMQF2ia189maXHkRrGh77sj7DNs
`protect END_PROTECTED
