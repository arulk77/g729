`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42H5bzKncf4I+vC5hIyHYZL79whSnlgRaDdtYklQGZmF
XR6tABrN0Zv2vw9YalirhXqaCfS/Bie+Afn14SO0wMvsMye6F+iSLt4ehRd5TbTG
sYheofX5253Qk4j4OLWAaX6ewfXEW5LCJj8APfX73bAckWd+zqw+RjH2feGiKqu/
6fw2AJ3chFpgnhwMsHmz/+QXF0uF0L71ZyXUsrn8LjkrP/iN0Eujbjkhn/ejplwF
fGpkOeVqLJ0nr4gQalEsek9UM4c0JHMtcATYW/RnogT7K9Dh8NB1vQMIQwFsMprb
JOUMK1/LFUlKkkouqy0WpcF2Z6/tvpBsk38XTiIZdXTPwMdErUK9n7jtrx1DYiQP
/TG2uemiTxl4MOKdvbeDLg==
`protect END_PROTECTED
