`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46GWjmRXe/MWdO//+MmMd1m5beiSDwslL7vE+OMrqBf6
CwoMQRR1XB7LHG1kW8cNOJN6nyWe6lm3VYhH6IbkgleQwPzVGHCgWpB88ANstq6o
GKB+yVw4949LiGmgFHZPmfjWn+rjxnrWhUZD6nEz+OkyQN9K0sFnYp4SAq+WjS6h
jGIse8RuBxWzni9KBsJEBnhQuKocOzNZCVwyvBU3gEpbkaxJjzAuqPO3gfOFVtfL
LTPCCZQv3/6tX8ow1Kh1aqWPD7jWrnMqIxuuRolw+3piJjZ+9PnQ9cUr277UDQpB
GsiRwfuG5crBhxYSOKCbBQ==
`protect END_PROTECTED
