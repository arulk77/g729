`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6u8vxV9AwG8NMRd+chpcM147H7Tg3eH9XOQ1lqA7Wowk6zYiFAEwwWWYqIqEtHSe
xM7lRdg6J6E2irtUOV1WGWwGweaVo7opm7ssi47q6RzApsjGwLa2aJlV3SE7aNir
IiABLh/5b4TvyPVif/3DiGpUqa3R8CQB0ggodryFuCIqaGdMwltQk6nBLr1q37CW
dZ9sdXpp6qso+s1sEBT7+IkNCS6OHj2860SjhXCcFkYivHIlihb6+SoSYKmkpTiH
A+L6t4YMVX3bvqIQxoKDwKn9qwMdSp+Bgn0r6Vm//xQeHHYBfg/I0ptyL6d2jHKO
hWgZeeqkgylST/B9fTKSCkwp5kpjDLlq7W3yLi/cyTRfGjsRCIrEnlQ5msNNhLs9
PdSQMDLxyvWLYD4fktMaRjkm+f6pR/TpgrKyk8ffOPzqBeYtnLvEF1Dk99U+qJMx
oY3iWVtY9SXCoDhJpGHnJnKca+k3bCGHLhiwJQhSEdW9M6bNo5d/ih9Opx/HsjOU
wJhy3B6QzSO2YfPbjlQAFUaYtO75DC8EJh9if45oYzbqFIvlC86t7dS5VSYZ1Dbu
lG6AxSVgc3ph9PYQlwHcvgYKn9WdHuYVgka+JC0cDJGBPSvYcilzrvwSyWqpNnSJ
mNJDffYR0otGc8uV7TTVW6O/YkhKe3F4e2Tmgb9aGDhhFSapZXuhPm1cNvgHZjhw
rdai8oE5h5dpnkrCwJ/dIXB0eD9vElx/pZImvL52jtDCd0Spq3bdUjahVhggbSbb
QMb05wjB1GjEVnrh35NnMMJwGk07xw8Jvf5Rrg77min0G6a9zihNwRfgBTPnJZHt
IFbg2q0S2+82/qRU4g9Nx77v4gaXgVe2nKOy/YEpi4I=
`protect END_PROTECTED
