`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveONLigS3V2HTf8883f5CTMKBQhr74dFafuShkJ/CZCGK
xlAnoiY43Tj4yA30lI2yx0FzeFiS8Ao9vTeImmnYAZYjXPveDDFqkUM6dLxPSiG+
m8K5mr+fcLkXDu09ps9zJ4vJY0+9sM9u+qsFEebtxP+T+DZljlKBbCfI8HbBersr
CEzuDVgHDpCvkKsv/yrpoDoYH7wTdBJsKEmREDbwbATYDZDbyZFO5YVXomLs0ESL
`protect END_PROTECTED
