`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wnVHZ+iRxi1quotedvYkSE2gohh2EFFmzI1ErmHS8eb
4j24mJK7T4dNtHBcVEUcNtXgWzu6qvWHELwQX/mSIvBRZZr8tMjkFmeKCR7S9bCw
Ua0yerjiLL62lnAAgDv/A5nlUmXCkwSSZyLmZ8MhWBwlD8zwaf7p9E3sRneURAHb
E7ym5Df9VlzAxIAfSFqAHoq2GhGi2CAZ3s1yZD9qXsGByt/l4dauptYgXERnWUbv
Ju3ANrNrbaxg6Q8qWVc0g4dbymc6eWkNOIISk4pimF8o+vVSVePEakxBmHMQGwK+
bnloXg0QsxRDBnPNct14i7Gn2/EqQ2SpBjJ/q5eEmz37uDEsaCgBhwWL0IAD8blF
QLN0EPciY4VtaV96Yp9aTT3fwGyWru3/xk3DpcgxVl7dTepjuR2X5bRFRGRgzPtU
vucEG7bSDjb9jTLDdCeDb4Rx3swcN2jaCXyTlGj4Q7bGW+yK1Aw6eW/PiVYKf8RR
Bju9BfQdYuXlqDsKeo2DcyM2z90hbMypJlMc0Q1XBss/JO/cmeIjXaMH2hIMRQcT
7v8QL7s2rUWFUfk2JYOFgc/qff9qksIF9VRYryIxMz3LKlcs0OFdyFLBvxt68HLb
`protect END_PROTECTED
