`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDcFa7UhTtm8JpXs0mzIwT+/5jwMB7+C/9ZiBAzP6Cj7
KV96j7sjfwupFDPx7Yy5aEeAKFeJio4jI09b4RLHJy9LT6SZrsIcvjM+UBlwkTEw
Aw3xStcRjqcEqPOjkNqTScusQx2ArkUtcyaa58C8k29wnftZACUvJg3pMHc2IuWb
epiYKeRbhBmKVCIQ2+LJhA==
`protect END_PROTECTED
