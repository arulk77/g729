`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDATQ3mJhww4LIL7uVz5N1m9l9n9HnzmQwCGhOezN14qzg
h++07NYtFrE8AqjLOSb3Au58LvlEa7d2Ls4+xYB0pUtddbNmG2AHg1cijgOH1sXd
ron6cU8r395QHhiO+T0FwTrKxptX13CDfo7qbUZCJS5i5uM6IGubEx3YutyV1MfT
Wp/YI6V8uiyZRBAmf7rduCyNcW+la8/mwQ/AuhA5yMYOgLt0vQrOv1kbpCsANPUi
RyecGhgNqcAGtC0SSEmcE/PFRFLyXm2KId704UdVFyiNpiEwu2KhVm6HsV4yTjKv
xwuu5hkWiGMxxh0TMIY2RlusPJxt+54mkGnCfL4Urs3t0oNp3w7ESuAF+tOs7MLi
qQ/DnC2aGndDTmcRj86mHs84cfo9/mGR7Wg+w5QK6JNqhPwjXeU0m1oydQqcvsuc
RViLa/NQBX4MK0c4O5EBmg17F2wE9SdxdCZmCpmu4Hl0aQrVfrymM4s+io3LgBl+
Vf6WqvwswYBIk/auDZ99YREDqm/xSrcVBC2IDXAw+5SKvv2oFmM6p5L0eFdsNnse
2vm+/1pfDIS7N+Q+iMb/v4Tue9Ni0yAIMQawnVMU/2GUNxewhwfCOZHvOWiAfk23
x189R1Qq3DYWDMZr+pjihg9+RdJdcPI6a3yMm6dj4LvWZA+36o+rChDrQ6yrp5/V
KQXIg4bKYMK/t7ZohHlqXwgc93dgdISNMFlo66UWALrAJ1M3mXDOA3fQv0RBvaun
jTiQj+gpzMHwwqEKDroS6Fh11SNt1KFvjGGoRBK0yCAVqi/cRs3YqRL+b1AqyTka
bFfsIxHmV/qgSD7X8cVk4WGjpGOGrRUp3QNynur18tliVuf39Ixe8Jtqdzury5Zk
ArGBuSALLNl7dkIdD6ainZCTMKXoOIdtNVF5cZcWqP8OLGmnLl/L+khHFxh4+j+r
9A2cGFweWwD0GK7gEZ8skZPWVrukPuICJp/o1BplDR1r8lxbQsx2EeO1iOL7ICRB
z7iB6iqMbrUv3bOJjHsAwvN9eKynY/Db1qF7R797IBZgyfW4qH4vANHiSuO/Vjj9
3AxbiiA7lekiR5W6yxeG2msUnm7FAQhamkVPF3SG2SFAJBR8U8kg5bYQSNhV/Hq5
`protect END_PROTECTED
