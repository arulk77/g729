`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+wF10l2PN9uSYF1dqrrbMwXF6rUU0+kD8bVZdesTwCg
aLbWLoy25nUU1AXdYH+PtzOgDaWUjvojeWp/weZ9DnvixxN2ezZorS9WW5ebAVza
MzC7Z4Kbyxdjg7dmeZjEQKHaJwdwqjNYmXT4d3i8CCvr1ChRsVIquQjCCPh3Ho7r
cHwU/LE5CdHXFJKHk84w/ceEWzizpRXpy2EVjTs2c6/0uhD4Dkf+s7pyHVilxmED
fTCzU7edHkF6ip/j4zHXjkH5YPKC1GWfe/IZbN2T/TznbiX3F8xvTWUAKhJqDtfg
KJOUqwJEFtrFJRh+7UbFxw7wLyqZeuMMY6YH2FWsL+JT5ysUBpOXngT23Jq/twL3
Z0WcaPA2o8CvKFTY8ecjZA==
`protect END_PROTECTED
