`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJW96zJtnaSNtN2FaV8LAaMtPpa3O8kO39BTROhU/GV4
s6bSdMq8kb/WF9AJat9Znwy+dFdTAnbSwNUDwfNS5SA+cNX7Vpx5S8KIo7cuz9Mi
8Rv1K4dKV4yBMO4RJFfgpVBPQkAGonQ/A6km34UyvEaQJiHmVKhl5/3hsEH4BmpV
yM4IsVdERZQn61bwyleWLQ==
`protect END_PROTECTED
