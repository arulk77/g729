`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP3g5v1jez9HkS2IjSGA5h+OM0Sy8ZCqMdyu5eSlaZc9
NsuRuFbf0rfD8L63oAKTzmk/u6e3daI2SyBo7KkwtQWzPUupXd3yyuWcjrCHNNH5
nOBaWIi2AYWkUVxbVe8UPV2i/koKeV2l40N6Bi+ZFB6X8vDfQx5YuMTgHXhMBNHe
mFFRCrtM1wkY9NjBl0LkjWDjRtUD0A4aoCsM3afHIOSdN0EoMxMactZW8jHa4tAh
QK8FnqgDV2SKCJcJs20ivF9GIkwVfSJNFS5t8NeUmBR96AF71En+/FGOsIEYZ0Ac
Ux/0P+4s+eFJFy1uYlaGKw==
`protect END_PROTECTED
