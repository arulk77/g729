`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJKAeN7Jo/UNUo4PJyNJVMHCt0aVSfs5H5OV1HXghUwB
iNppDDiBpCPkEIjs3o51oqk8ZoyZoJ1KU+/hDO3NiShnjbIq61ONBVvRT07fzVrn
EEr8ZWJVP/59y873+tjJ2YfZb5N0E2hUaVZiDPOzBtUPAUnyQZacOUTPj6b8f3VH
15i49k86iQW/jlTYDynH+dQmbbpYfv5L2JLIT0biZ0kxa7aEDn/7Zdanx5JLRzEB
BddD32HHrLbej6qY1UazFzChrqyRQG/b3vohoSJUH3fh2ljqmHIeDymcfxIKVWOp
Z57Jg2dB3LMlPkq1ElFEdywwWuhJPKiA4nD4yTqEr94oFsQ4P0oxIrmqPmCV20Kl
WVlop12/47gJevQCllvnow==
`protect END_PROTECTED
