`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GnozPa0dOHRBcNIaQlRN3ItHtiS+kqcn2SHvEfIF337xzI+LmrYuwUJ8jO7w1GGm
pxoun6X2BPetWdC9JiccZ3TP4w+ynT22OwXEqzUdPTe9jK27+yJXKzlS7h5I3gUY
ChvQAFDImNF41pZ81SpihM1T23XV5lZ+WZJTQYUZL5JtW5n2922iZffqPlBw83vX
OnZJLgVkns0yQhdz2R8HwiO7bX1e20EwwxmVQM1g8mklXy19xtLjf0xTvHv2IhLK
036Ze+ELGNuEuJD+j98NkYchshUAJUW3+fLUbzXCPUKQph3VDYj4kY+OxW25iz1P
R/zQp7Q7BhD/DsymM1QdvypWz1fU8kkxwF0vhsw5RlYEUGcWwFYlALv69nn0gHzZ
DDhEVjaFbouq6t/jmYLTXiDx4OPSC+0uy6tM8aAVCNOKWcGNt/8SsicBQ/1uRXqi
hP2OD7GI0ZYgExL/bFGi3px2e+qzbMvuQMG5seTj2SjwKjd74xd3zzpmeJHcDd73
cFW5LgKMSELfj/5m/tK5W8QMBsIiWtOqWmoVOoCfhEmLAhia+Unc2Or3a6qOXNeB
WWG5XYxZD6GHFcPCVwtS2U50Jd+Nz1MMFwXEzcyH02z2KWkk+t8DMJvUc3AuuNiH
KGO5FtU6KzRmkgeNq45P0+JfppNW0Xh8q5HPb68OoGBL645fT89fuOS9yVYJHN1G
WqK8FhimQYeJi8yTk54GAvh9sU2r3Z1cjsd7uqJAcQZ0UVJuoags0rolOOxFFXH4
0LHEsTwevxy5/40SVg9dsskBnebk1sz25PUdFzqgOeH28La2I5j/zxmBkt87Ou6r
s+yuWomvXzYb1vTUW/f3Dv7oHSHLkv9ia879fpf9ZjXyADStOMZ6WNd8+tcB2u6p
qdPqk42NJt8a5pBBCVdKUJOlhQSUQRbDZpZ1tX9ZR6cp2F6K5et40LALdKEdyf2y
VMwtTKSZfwU6uFPUcNaoU81MrPw/+onSKhPdagrrKtiutfJc7lJI4IbO0AaXfqpo
0JLXutQSVrXooij5GR7COZIbMLJVZbqkpmAj67UiNnJxA3s2i4yr8ecQM5Qi/+e3
c/Ae3Z11eC22DEt8W5zIaRCNron8qFyynZYWRJbzj7ga45js9+xjW5nzxM5iQr2m
HaLt5NtBqBCmPadb7k7WWlafM31SyDCq1z+j2YxUYCKHHhK6FURnXhkmHGPDJC3T
z2qbmSKhn2eEUKqqJKpQJFC6+KpvEtnc+6ziPk8OTTx9zP697CinrrDMSbFLZjg4
SMubtleW/uYW939pLzdZbp7MJQpAPn1l6c2m/KMY7Epd/kS6wBVxkoRd0Jx3lXVr
CI0drCCVzONF+Yw3A4v+Sv5Wf5zLFkjOFZ3zdNKCDEQrXnOSZ0XR+FrqUKhTR5Ma
7n+p1I+/bIgCIFDqneZHgyl3U8KKJcuiTc7J6Boa9ASdfzvGf5cjIkZr957IxMmC
JBN7GmSrNAww0y5Um7Z42uN73B6xosj4yZ4PohXf9pUosrrWZEof3cWq+AJrYozp
K4UpWDcpINSB3KPn92wR4At3bdwLzpNq2G6Ves9w9sTjINDtzFYkcAf1Naiz/Mq2
iOdAS5Uk0D/gfSHwcNnPl141z9W0SHvc55D6VNPyegRR2hRp1Q+4U+wsAp4h/dEQ
xwsABnJYBakHDdMrW39uhMJ3JXRMGMRyu3Yj+TA9Kh5HWUwyxpX3WznBr9oixsMj
OEPW0uHZoPE3sFu2REl9C1qEMncoaOusSaGLjh37de+vJTAhnx4yDU5jJ/vFpB59
DMNqe+POpS2zgEYMgUPFWc0pc/almKkRpRkzTKJziuA8lp6IR8s5bn8tFSxERe1e
RFgvz7tTomgIHgavkjAmQIlQ4miXRJyla9u+nCVyLxh2O/D842gJhdUo4wl0UyEm
fh281zadh96xmJHbbVpUrzSf1scy6vjP+CF2ijSxsLhFLpuih8G7KeHOM6jjkkSU
VXdu7VzzlEL6kDiXQt6Xr2VTiIKK6KX9vyHbUtLyIX+NpA3p08dKPh4ysGYs2IqE
3baD4SW77s0vKdbSnqjpfwBWXVPWob3MQDJkk7JELRMPd+hMzQlU3NcXIcE+8USp
rPBE1RDLdS/WmXBUaDvJOEsrrqGQsbDKyQ5fECiizZ4orKaFQjjmhRQslkTCf/6q
rXLtLB1XIhzeHqQXAZE6GUHJhJP5yyzvvfX5LRK0FKCj9/6kAJmIo9bBI5pCQUF/
sQIwnJ1eBZGpYc+H0VFBmWSg4SSrhiUxs3RXqDrDG+Rxh1xli7twexlsyDZceUHe
lknLXdemhKh2B5vEZFVwSq769M4Zoyz46LA7S/MnEZoWdRMbC+V6OSTajj3+zVQ/
jjdXTpDASR3RHjVyAbQUHui9UyYOMZJxlgQelgy3FqZMY/l1J37GQj6Hc5wK6ds9
tbzrPZGiPyb3i4LlVEInnVoj7gUbSZ3T5C3HeIfbmCwKZAHu9nbwL9wRNRo/W1ux
Aab+CuQhq5x0lTiEApl2+f02Rr8zUmjlUbN7rg6eXns1Yp9xDmlZYFfRi50+2WpG
wfHegvjW8AEPSFnyEwvM6NDVIYM4uXF3kVoPZm4c7+qwddtVL47lmk2IipAikyVx
PlVC5ooyrGgQZ9+bNwVO7AeZhJH036VZMFBO9EIy1pe8vjcMTgGJtUbfHtQ6/TPj
RBCV+I8eT6gDIaUTHim1LJXM5uMmGTiHuGYyY49uyFCXEAAw8uDh/axbsoHZb3bb
LdkQqFyDCTSQiRlFaiAz+gDCakZkIeLUOeGB22FfbEAe/8DD1b09R7eRaDCyYcR2
EjJIdesRt+kntjy9YmI6ZlDk3t0FK8Fhqd9t0nrVXRkS26+gec653Y+dpDZkhTMK
9HcXzVwHunidBWqMF4T3sFUeUxjzfEfuEXIQWhachCXqsdqiPhOpUR4ahsWHy6v2
MvXVRymBBIPIz38lN3g2/6QECkmJOzVeAqhuqO1lccqjIV7cEXRKHlwaJqo7dCqT
7uXvuTa6HdgBPhVr15i6yKga1h/2ewIOQjsZMCsHBAYc/aZp4zxOd9kxLuWgMY4c
ivk4wymlCRD4qe3Xl24lgu9Lthlxgoi3NPbMUlBwcpsN3hVhW8+VuvJ4pyq7RTzE
GKEe2VcyKkhXR93mm4+wMY/kiqfFrEqnZ+bJ6EkNudlSYpRHdObVfrRFYm4sPQ8U
lpoJ8ZIa7kOqtdYxDxZwLGre9ATph58f5N6wK5iwXWmE6bWTV/HzhWBb1ErmuSgr
Y9xlyJSeI9AAfr6CI5dCgYKUbqBEcV9uuoDWduOO2e8EhLJrCdtEXlT3OAt8f/we
50Sbnar7gRQX+MVQ0fpSICxzTfICa6cm2DURejAKEn6QLROMJ4FQ+TMutawlICh2
1w+c5PuXJYHB/OzNWe5OYHEYhGEcc8i+oSqzo7z5rlSJdXbcrtUod2vtwdzYdd6Q
c1HwrEKRP5SfbvOQ0DDaw9sVDXE7HXIyD1MKRsJOYtIDz5zwmcc+ybX9DBOMwiMx
1IbPhvsnoQhapN16VknU65A78saRT0n4zJf+HDmDtapdQu2YZvMeVd93c466N7Zv
op6KbQgw8mqnnPTMJDhXL18SnJHsrQjY6sCIupDetBVIT8QYyYKCXHJj4GG3bqZi
Z4aFuYclPVzMjaB/JogyK/sqCelv8j6TwKsT3o2+tl+ZUIB4rzd7saZRgaf1rSQl
wJE0+Xhsq6+/ihcOizT1OsSGN/von5HsxuvjeT1MbWOiqQt1s9V4pljJWEpTfoly
i+u+ksQIjuAKoLOOZuzrgcHtq2Ss3+IaRoeu93IbPDcT6Rb2APaJg/mu56VvzyJ2
fx/x2Ux+mjvVAFpC7v8v15WUQB8V8L/4izQLjLFhSp4rT90u57O/rfEw7ACfOdFc
Bcbd8l8BaYLjbqn1UNocjUaQQu9J5YrjECW9XU8ytizWURiKMoz0gLx0bwZpdJIt
cVHDAMqaHRWFoUgLT99MWNTI7pivrTW+unt1/CM+YZwqSbyiFwGzHORpn9QWcvMW
jnH8tOJcY/Dg7i+xOWOx6NrAZ0GnQYmGoKfu7xr96nLz8Hcz4WLg+eP5aeGaKKH+
4Rzty4DVYssrqV2eRQXtJfTWRlBWM1nQnrfJoQpBvBe+WJ7n0mte+ylk0LP9HPtG
y13sMD8Q/ysCmUhrmuioN6HTiAbOzt0TF43fqC4PiVaXCSentZ/tIiixJDBA2aoE
A5LcyIF2a++j49t2rGPWE8r4KivRX5KWpfg+wfVFHHXQdCPQob/G16/596WRz/DR
+dzSuZTvYv6sRY2kP6PWRKYqAkiWhJP9c962nFKayNlB9dU1VfoYSh7Icq9zuCwt
3evSrO8r9LiSl++yTRXyIbJTJAu/TUCNQ7E8YFFwzFV/e605v60U8dT2v2gBlKyG
TxJVloBazcGbLUZo5WnXsOW9exodr5F1krou09eqf9AcPoULWjaa4vctyNv7+Dms
LkXNh+YKsDgEU/UHsufZG3/br+PR0qork0fdczCc/7nHG+yVst5bEe0NDdKuwSmX
ZRlxVSmySOjssuPPlUJWF5L0nbixA2HoLexvcL+k52jjwq/5QxorfKdjKCAAd/rv
L6WYx9Wdd5Hs9ZRKypjXbOguJhrwyTucSCQj41xHWPkpts9MkAFLD2lG83Bil6mb
fJOvFXfThI/SDYUivw7/U2bc+zE/glOiS0lnf8aLmh7ok2scpNfxu+pcJRa0gZMA
IX1ZIB5Z8xyHesYI6p4iNnDstmHQsPR+91BlV7LFo7NDP4P6cGJwrAIiCjg7PXZk
ok0pCnO9TUNsmtnmxKOEv8BF7l6iRmziJia4s8mebjE=
`protect END_PROTECTED
