`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RY/+Rf2AZ0W+MdVJqdhaJxCSWqN2m/+sgeZW3x5nup3ojcvHGfb/99eUd3TXxJcS
1cfBCDhHUsqZTKyg0/jkze4TnB1Yatu74d4PuY+2YEl7ZBI5c+7WH7tYQhov2a9d
KoCzTPutMj9osbz5XI6Kjua9RB3u1Hmo6nyyWaMeCGGFpYZn6Usj6QkYSn157m1l
naZpHOCKF07IylRPv3yIUTG4sM6srIgVDFerx7vbFXxEo2f16PnE48yJAzgf845f
WCKF01Kr7rMWyL+toED6IkOF0x5uyH12sTww6OBZVP4Dr3XJv+BcCa3YaNsSEET5
KTqd1mrwR2JpYNA+HfhDPqrYoPjMSS7yqgFbaTzzrw3UYQAjZTA/L0qzxBXDXrzz
x/0soti/w3HiQ0vXJNQyHJsj7+jz6cKeJmXGAUsFxHGWfz35l/8qQ9L2NJLa2AZB
XQB6RdKVRAnKwN5V5CiOmeWw8TFO7JfPofy+zf+sZAjlAoeYYlnO7RN3XHGhHdOa
VzceWcJ5sOv1eUXlmTQ1qJ14nc2zmQeHIWx7q//QWCU9g5XOKZaxVPTN/fB3Hb3A
bxdgdS2ShNb/Q1CnFsXCsS1czaujeTx/L1DOCru69dY=
`protect END_PROTECTED
