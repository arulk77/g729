`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMN57yQVDrMdt+V1UJGcHDaPeXrWlgEGivnffzeROVLK
b/NbtDkeXO9WBiCGPuEBkBWqv+Mky3AMx6ZwEW2UF1X98RSnD/LxMy+OU/Ujg8ig
OMtCy/T/D7Q+LLFTM+vJYUCpQFN06Sq1LmUV5Cld3JiyIEmxYoNqnw4uQDOlOYIV
3ph2U2bJ3hykCR8+HXErUQ==
`protect END_PROTECTED
