`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePkjr6QNsCQc+IaKW2HEatpc9Y18ffbFR4t4Ggb+ycOg
taLQPkE6Qcb7lUv9RX9ojFuSE175n+VtH16VGmcEVwvuI5Rruiz0TH5/hAlTWz9p
h+BLpUHJdpUMGk2Lh9V2vRnu7LrEtFW/c5W/kOGkCs73wrH8i9INOgZ0Zw5x2hzx
lgrtwqCpIZp/PRJU3OrB3ksSYP4IbA/qZA0ThwYx8EizPvtzyAdjXElTeNmxtSD6
x1gggNlss0PttlZuF3ANj6dZ/ukSTku9QJfoLlpFrpmnDUxw7/TKvzToY0wyUx9B
GtuUD7BvHs1AqhjapdEBvebGqFl2JSjuzIE6GDWbZ4a2eNdpxPGp6XZLm3AmcHQJ
HTqiSztezrQm94qrPKAlo5Akk8m/+bZ8EpIChPFRLrSne8QcfJv1Wnco/V82lADG
2DlSqSpr0XU/6NcTcTs+8s+F8cFLBseYPPu/Ej7uJQ0vDP7wGeTEtk5S9IgR4fso
1J+z1lyVH0JaDQ8jdzf8aQ==
`protect END_PROTECTED
