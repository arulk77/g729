`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
HtIqHOeaIpJ46WGlN8M1OEtCORtcKK8AVjSJD5W5xcCb1gdaLZk69TjZ0inxK6Rx
OrlVpq2FynB9kI/PLz7TDDs8saspjG/mx/RO9yHGbvIEFN6YgCr3HHEpvHw2g/oK
hLtxGnNQqWbd9UbkOUvwx/HbVDqG8K1USdQ3W61wuLm+F9xgsaVjjHnaNrEAA0Vc
oO6LVth2SYcQXCM5jllTbKzHPW0wreXvqRLEU369Dj59OX0n0fkj47Rjk6kyz0MS
jZYFmeO9DMSFNw6mRWP0YJ82mzDoVWSobg+MuSOQVei7z30d2P04rBxFcG5ZfdEM
UsbqvpjXv3WoKDa6FRqd2xxkDhwv7jCceeMm+4GiEXVmRBbzL+Qz7x1zQGOyDoqj
R15ZQWCwlIIq72CDpfrARCW4mXM48R5X3K3GfpOZTNJoCxWZUflreaEyHyxoc7Vq
/pslWkQY6RYjPfNs/8hIOKRpbZr9393tsiJQBQ9OOCuFIPP9GHzILefuFBUshfuW
Va/JLTgTobKMEb5wSYweT9QZE8P2VjJar2JY/rQHD2H44avzBClL6Jp5PoH02ley
COoT9pMjPG099bSSdlqi+WTbbuzIaR5heHKUdtdhqBLZ/AFWMkkqpI1YK2AgOu0a
kr6KOGnszzKBqNg0+oqBDMGQ6Avk7mcl5n8ZxFTFcK+UmVn+tuDvNjfyKl08PTgU
O3OBaoEbFXZG5fmF1sqJRnpANCy4gWhd+Mr48oy0O/cH4U3CaxVKSnouv4bodEUR
g0c0iTK6rdxEqGNOqtd/sVQeJg8UZHjcETLjAY2aN46r4SHEXec5UhHufzrHAc4h
LwaBrkvjOOG02FUMnCgPIpNDTbiQfZDmpU0lfDMLlTJKNZd9akYRYJgkxWYeLz1H
TqeS2vsxdKqtc4tDgHeu+UjweSl5kg0LKODpm5PfclWBwR2rW9qTt8wr3O9O7Ba/
B93vxR3TM//vU4bP2/zePks6zNHRReYq8N6AHuAVYLF2mn0ZMvLSOvYmPh+VznAd
1a9zqWu8dpi5kWOGmpONpx12EaufZFcz73SpLGsvR64Lh8vyvH513bFp4Rijg2ZY
zXqW41UnQ8izsx/H8AG9QNlk4c/wLwnUM3ooerUjDdoDIciYJDHtMnv208AE9r0r
lZGTx+MPyHxbpSqSFGu/z06ZJ20rdE5yjeweRj0NoYY0sl4ktSTjor+jCwDWq6Fc
u2luYo4+fY815G+FdW7v/qYMYBKpDJWHI5RqR3sBXqTjijwoySg0eNUq0tzCfSKR
ZQgTNyZjsuWDDueg4hoqs1me1Eg4WKuNFPKXkmxOYqnmy2Axz4QCDfnrPwbpaJ2L
dcemaXFvRV73HgnIqMpIb46xPkAmYFxsEH9Bo/eLDn8ph1Oz/1AxqDpCOU8RMEhf
p/R7crV0gVvhKKvG5xfKdYg8RdGZbQ6lh9/tACxF+fms6CPd6ibkWTnMPionk0a6
s/3Nt4PwTRaJf6pOg/YxbiO9BEped2hb2SDm03bJxivbiWHvhLtAFnB0GGaSiQzK
yvvPIou24WJ54U/ZR0Droz503pJqh87X3UwhD3glaEXx6hNyt9J9AHY3smp0ixrw
lmchJTkIOUE1KKQwXBu/i+95n0okCF9SaRQ71Wvby2Y1BXtxb7YRz/3nkatcvJtK
9CEdfvKNJDM5OnEKB0nE1Xx5NQpl+09O6aHGiWNBvzP2WMWV/VkfMch7qDCwewC0
C+92mTlf71P7zHZCSorJNi+PYRq0uYQMyYHWBH9AqxlR0IdRSDixy3q6vECXVxHb
/PklLR9mComVET9Vc+DFIQtHFscCwzm18X9ZD3K5gWE=
`protect END_PROTECTED
