`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41978GXfBnazAzHzovRRbWMPrpyxtE8OG9o9gdGVNcoh
itesz8mQXmGs4tbOqoU3NnTq2Qkh8z/EaJ+iLQVZduR3Rlp1Ssv6e2o3FgljvPCN
/eP3SVfGzOmxkJ2f2M6qA4xEv03glF+W9/AWxxIsY4kCiOGeGsgOcvJCwG49tYqy
5xfTZIJSvLWY+3vx4S13GpcBQx9VpfL3q73ZniSfejOeRdr4hxZDuEfCH/Egyq34
pYkrTLMURA++GQTELfCAhASaXcELGEjPTEfzwlal6d97pf1lx3fwbRCgGw//Na12
rE9IywCvYL5J00cJYjiBeA==
`protect END_PROTECTED
