`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePlZr5BcU/XbzTMe6WdOwa1qanw5Y7ZKV7oYt/GEsXzn
YmJaRYeWMa7Kz85Bd5+aYFaTElQ+kzY19+LrWplDONtQja44lXIEQfXG9cRBu7QS
jC5bhwsrwJhsCCisT/pACz0rRHb09s98Q3OUYtfZ6WIOZNmd73DjiZ3H6AfyzVV4
pIJ8C3sZmk4OE+DJNXCdP8w5pRWi01a1O9hhoaWG95k6hgh3d0wbWbKYLmNigIxQ
Y9kqBB8DXx5MmIkqNJtFkVG+023o+p6Kied/dVMBipUAcrYimmdpqf+/EeGw4ZEX
c7MyNGW/7338LsuYcV622vhnfM8pnJ77BYO8ku8TuwWfIM9OduyDgMGJ6g8vZKkL
5rR3zQJf5vk5voV3BMbPCgJ7J2KacQpwhwkW5Oi6S8nZJ8OMpqK3niFGkp2v5BxV
d50FlZC1I854OuTE0AwWTzA9yzDiq/Bq+pifZXpRD24eYUlu48SvvnVLCcU/RVzm
uosviZ0yuMEB6vxx5Jjsgs5aBFgBwjJSY8x0LTCPX2A5ZwMXu5BbSw++pnttHPER
48hMkvmwAaLBrvZbScO9Mpto3n3KBUqOJZ09bXmWH70Ant1QjhOm69YK5/yUoBN+
PAGlJSSbRIHsTv1NAvoEDdoEuZQu3jZomUoZDDgM1CtfdTntTczU9tP1dvSTmAiQ
LNVyhIhM6mHijfEDa8dJElO5YuES5QYyF9khS7kYnWZaBnPo9qiIXOa55GFB7zwW
vERK7fysHUjejmtql0CXVTpskuCN8f2hJ1oL47+cUZ7lzIdTWD8uzdcvEKBxYvFy
uurOqBgLr3k3PGdBDo0ijjLq8Db6mY6GgVbABFkXM+U=
`protect END_PROTECTED
