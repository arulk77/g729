`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePklW2jT3V4qaHbc8d8Tw0d8vnEPbOcy+JYq/qtxC9RZ
7c5/5PH3bhZ6pIvgriLFb7a7k6Bd1j+sJ6vdBAIlx3oihUhHMKnaTlm8WqeQDgvi
ih0maOWzFyEyo64aUHeBZsRpxkLX3GS7hsiPCU2ERgMFu8T9MU3jmJwT2r7i2bq5
Elsl4RyCei2a9UPHbtGlruvVSIwzBi6SAqNJVGGh55imZyxxtl08XHU10YaNnSPy
`protect END_PROTECTED
