`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLBOIEnzZlSGizhPMR98roFNbaDl1+JVYLia8ys0Qo+V
qQnBhzCIotInLoeOCcs2jkk/FQF/JaG5Hg0iFx3NcAQNCTkIsUtitgT2jGBsupsk
TFpgu2oOpnKwWrKtj6f1PnY1+Cwud8CsfmzO5UaV5dv77LLNCziSKMHZzWEC08pm
gbTdAz0tvU3QpvAEkU0TD0dIspdMUJV2riNp6wYwMK4OVFqq0GdHfreCeYKFwOAH
z9GtJP6iWj8i1z8GYRcash/soHpOtWTWVPb77y9WaWTXNTbm+QKfD6eIrDa2E7x+
sFKaOGrP+4RNwxM4s0gQ2Suz3mMfCV1QBj+RzOZ1dfc3R/i0HTE8I5kZmLAuxeYK
0Dln3Gub0PzxsA0k2JbH/P22oWWrNFJUZ/D4v3stoLXX/fcI4I2k7szNl+CrbhVc
a9BlsFp30QFt0lj3DS9A21HVdcHJbkPc0nw7N0FcVePSmpWMa9SbKz3d4S3fLWPk
+GB0C4IFEDzrH8wHQ8gZV7W0XRS4Xt2hq84DAQ0Q2BdXUdsG2q2OBO1j6GyR9zF8
`protect END_PROTECTED
