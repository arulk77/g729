`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kfggrtX2fdaKRFdv0h6+/JhDCVd59X3SEXrkxD81Un8gM6qTBmfKAqd0NageIBmU
Ezb1lppz29aLSKT804nYp31KomChPSpbbwUVfA3yPMgWyXAvep+pzb042ZX0IkE5
a+5jB2EA+lczI5m6qV16gblGkPjegd7CMTQNmZOjCUJnkue6JNuDsmuN12xqbZPp
QnNpeigWWIPQ+vIUROkgUOd32AJf13XY4xoVD8BONHImNZn5jJrDwUzp2yIwTn9P
blqnBNbkpEHAH/T1YoCir5uryx35DGsV3eXbtxH0Pko=
`protect END_PROTECTED
