`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0UIQ6cMp87wJIP3pVJWYmMo3EbUB7xkvlR8Y+JuDzB/
fwEAjsFXIbv7SxVehvtnnnh4TvP3Fx4KCBtdAAQNU/0KuL0SgmN8LXUzhbnybyfg
k0vqlGddxLgvGRX8mL/PJ1LZaThQCdQjuoCt4YUaE7zie70W9g1EJs0eEOOklHvy
Snhd8M0QqQUuAo6DSoIY5nu3jS+jq9I+icHbOD+E494rvMLv1AYfEJYV/p8/PhNs
VKDECqEOd5PEk+/8lzILbuyGvQyKhdH78B+wAVmiKbHgnOTUsYSqNQQA5YsOJa8f
Nui98cxY7ulXMcEDhuj4zUlqxOUlqh3Kq0fMx3o33MEM4od1o2oXCeulNbedjrhn
OoS43QLsfPqOJfD1XT1svQP3ng5K4pZcI8euR1FSoI/Jpiad5toaMaqxjFR1YFQg
nh9TPuQeVUA2hpDMcs+BJkz5eotBvLU6lQWhfrPNp8SU/M2fSMAdTmLYYt5wMPtl
6IOxtR62igU/xo3fsqx0V7Ku3e1KQJgaK93UM68KqhuPXtKlXs5b1rpBbxVBcrsc
pCgfGdMX53EftUwrN52fmH7K3uuWvDsQKmuAptittsH4xOyLlfUM3zJgT1KJ/j3/
eJYoAbJ5Gz0snojOcMSEo1Ec2HiqclTRKRBsf1XN2B+T505NWVISbOJ5r0Ufqv4f
sJQDiibui5TGW5JU5qz58eLbsJeZc203wcMA4vRfhT9Fa7/LHNrQZvFh7snNUudI
2u2CdQivFn1JCIBQ4TPJKB96VsvIbLymBeMm+tIHzLe948CWtmWun5bAdDUteNQw
tLzJwy2Ksi4o0vW6iXUt/kvqUIiHoVLmH9V1rNdfEZkhfC5D05JTJeS2Mf0iLF3e
sYjJsz3Zlisf93maSKZS1gGSBtFZFr+Hr8cTX64/TKFuNx4uGRuztRK9Ba1p5Cec
8X/vvKHPQjVbJM5/FcuvXWHsJzLQNgEksrI3vw9WavO6+Dblb8IIep3ZXbbUd1Do
IwUQKOtSnfQGj55V0EUlyvBlxlsumDc6BmHsNfxJuG6Cwr5T/KTqwmDlsWZb317j
MB6Gi2mjg7okjtD6RcV3CjzMkyoJo5oA9VQo9Au4vMfNoNprHnYAIDuUMStIRCe0
FZ707AlOFbfKWuyZ3mJShJlskUHxbV5MgLXw1woQ7R6k5zOSfjUqCvakxml2x17Q
DyuWzQhX6qiL5GxLHWFHf8yXQvKYuMmJw1IAJ1EVRoXrIPnqFQ/cf2QcdoKXiptw
5zB79xLm8zEqs5sjT/8QNHVNPQDQ7BAHJL7SVoctQh6v5v91ZL7V2UmeZbzfGQXP
RjJGpnBh/brpkq6kX+5J8Sr+Q/sSFtyrwrqZHm7C8Czs2p6YXozjV/enmXaMVG/U
ubNZly3rLMx8X9jyUikl9G4oGohYR2UmBZyW90YPHDeutJjGeVuj+RI91WmDJW05
3AKWnpAy2YLNTbJDseWrt/HkvtaSWPShtcTi7hmfQbIzqgQaa/1AVW0g1ohyLd5Z
4/loTvZYj9fbUSABmp0NWgyc/K9l4Vnj8/WGZeDIi+CRXH43NUPhr2WP8NLcn53r
2uVhkA0ytJs685c83+GutoQl97dJ6z1ul7ZmDzh9C/o9o+R+UaRFOYSwu8TN5qNE
BY/tg/FB+PNk4FgskxYMcHnzyujv/smwpn5BIXen3AXDfDmTzRBsyMjUjMcO9xVl
13AwkuBAUPvVj3RBVjzlTx1/trNh5jm+3Rj7U5V+j/WMdFc274GEDk4kkF6bNr9y
E9VD+XggO7AhqYosExSRh7ZnSDR0P+3cpOyGd+w7z5IbRloXnJ5ArvZFlKMec9RC
8htyGa9N2A4fgpZQdtTlz3tZsLHFk/mabcTKHDZVvphDOREyHcPYhmtpOfDGzi1F
Pe8/rdqmQKfMysqlsfEzI0/jZ0vhrRvaLN3gLBH7uQQnQ6rOoWN6CpwnRtI/kJaY
E2/O9rT0AASu7mx+cqlnaYevlyPylku5Bqdl66lB/2lEyk/r6ObWOPXt6IovcrN6
gMZgiPawbPMobqlVG4IY428gyaeQlNuG/v6B5ec0QpK1bPkELkXQrzKOc0DUvcMH
eGZ0U/icxd3S5o8DSHU0XYQri6cGybQWrfv9pUB4z33lH5BfJUa+yjcftppWx8kA
JzujU6SXaFt2AOwywZGi66ZVeEL3qHCWeSxoKi0shKLkoSmc4eHcx0NCzU2Iysxk
amtwj3qPj5uwnpz4AXC516eixQfXEi1IRLTvXkYjaQDWIchY3z253rNEPlnUw1Ol
EXbD4VYdLsiagtUforjW1VfX6kR3Vbg3sR9qOoTL+ykGTR3FhoqyR8ckvLiV2np7
EDj0SM0rGPQ20QEVh38AFtSa+hwO0a1By+riLa6RH5XRFziSOj9uzUi0Qt6B2uBo
1g3CDBzdpioBDO7Db3mLYvyTziQXavDgAfBlU64V1F8xREJbZwLKbymCJbyTsjrI
ot4VRcIHXHy3AYfYSt1E7QxiSx6Rv3KRhDPD3hTOazqKplzPE/3fmyayljZ2t0Ml
6VscAShF89FCHMPvhpeXOpntgu75ryKctfUfWWocP3zL8eO2vj37gOvUmecy/g8V
NXjVd/JM4aQFqE0/0Dbn6zRy3nowuxs3HgfuTyec0awKpyvjj1nIgTYWZtwYvAAz
YK/Ux6OPSlVM13xiZMNyOLMox+udeP7lN6Fj31c/4VAPx+EZ/AnUsWRGvurQjOx2
O28GKfs90w66ne5pwpXKKVuVVpD+VnWcq16W8g0kKvKRldIrelf1BVIYe5wm/4qG
o4nxF7dqJvNDdxoRVgUxZCYZuD9uRsqs6BM5NOOJ7ld/LFI6NbjiyyMhllSWJbEV
PH5g/Jt7FZJj7z6DyoG58wdoq/0PlttvFwm+DhgDUx/RSddT3PqUmZgbkfF0R3yT
lsHia3NpGgFIpnVx3haElZBqDsKcBOvV4KEj7sfskpl0bshImsAIAVPh+2RpSW91
uH6vr2au8T41S0z9h4VzL+drg3vTFxJp0sLSgxtTMkdAT2ek9DALzVAXvlbaAefw
l7olhSMUkbNkz95TD7cG7iJ1BLRE52aRarkwlxxmj+tUPmDz+XNU0EQKzxwmFNdi
B8CBv9RZW1L113lp5AzpZWrx/NeMeHBz/4HRL2vlqOFf2eQwjB+sPtqxCP5IfSqN
UjUo+OfIHVHKcDtWlsLLloNlVUPIuSIbvEthqy6/eAtguy147Lf/9JnrfkBqd/g9
2zV17oujvwxSqWsDoQiWd8NOCq1voQ8mbqKC+pTd/69tqBHrZvsvKayRag+08b5U
nurY+wqKGhr2QhZ4nvKJksCjsNGL0AeO5+syBWgNKSjrkcDbT3RT8s8QKvRP68M/
kDfTp8zXLcFramGOqZa+R9iQanlbjNkPE+q+XH1MNO+y/defDpro40ThtQq66kWQ
5smFEysBq47urTf/NTE4Ee2FvbEsCxADRet/DXS2SK7SuTZE9DWAhfjx5NmN/28o
LkVZYZaRSGoc8A+PszVYlDfd1yQVddH0ZiS+Fv49g9pkLBcaAqWSF9WnJ5SloCYV
WFjnY1IfdAvA+r+nDGP90Fqqj9fAG/5ghzw1UjRn98nDk3qCRir2e8+2fn8U7Ssr
xXPwmNrtQtFOxCccpkekJMZvhkTWqhc+639jN2IWOBnZFAy/6KxDfVNviyRdp5Xv
Vr2/oTx+bdVv/7TXY6eIc0HFh6CzfeKN8sKG54cGDsLHY0Q6ql4EUGRVs9GaYk0n
uxfUACSUM/m1HpisCWADoMM/xJnMUkwnLvFI3Q5Lh7dEYen+Ul0EZC2JyBuJjc4d
PzPlxmWl0UeY0q6GMXZTp0jsa7ZMTgQLrie6zuDXQita6VpckpFeYCnUzxo+CIA9
C6fz1voNH2WpoN3+W5XhkhwiE3ZfhovMCDEUiXyZlrGaSfNPuOa5eVHlk0YhP26v
JdfLhg0qef7M+Z2CA3k5hOGt4yjcO/5NAJzYM7Ql313YwANjxyvMQpHc5IPJdTAu
tnqHWV8CMLfg4FEsM/eXzlHpE01Lq3HiXj5vUOzqTsvkA91TuSmx+fjcKKulKn5+
I6/yhpDuTwOYFoiY0UY5nHA5Df5Tm5BoJHXxTJV8K2WEFl5nLNJX4tjIuntHfdG+
t4GjgMWVIwLNnHboQ0/tJKcvNMuPhroh3EwKwQw4eT1kWY6pt712CD/XnZBE38Pk
7lY8NiqdW2bx20rUxT6q3+6X9qSBi+4qkl84V7TQnZkpnz38QcC0bFwxZb7WOqm3
pVKHXNmLJyq0Lr8qNhLJ3hDGHwvzPqickFRrIvVYF4dbKzq/E0JV+0PBS2qFmcSc
a07dP9btQFZSxUPT0VFFP4oXmgaiLUcPFTA7uXFk/jouUKPh+rvi5JHOuUwImKYk
0Lbr3QQiZOtkqScfeqUJYiBpcNbKjrUlWQcLPtZVN7J/s44W8vfBqtuFOYtRNBja
`protect END_PROTECTED
