`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePfG4LYuBIWaSIho/4zYKsf6MURdBqo1mFD9Xkm7peBO
Q3CKJgU2G5M5CQcYoLHhgUw/gWwZy/5vIk1aZpI3O/tbIGu47/4ZtHz2huY6Wwgu
yovRV89BytcWKg6szOXNqzQU09SENzcxNN0IHRS8au8HmHuoGhjKFI/fQmu6WaeG
+3Fwy+glj6xBlCylcYHCc/OCwUtCy8R5h9MFyVuYEb/WWlRuzTX/zc1zywys3Mgm
iApK7LMCkEu8z2SZ2Zb+fPa/Cgv4Sl495yEjv7BGMwmasAG6w+l9YaQ/AJo6I9AT
pbyJhPQoGi3D9Io6YfYCcw==
`protect END_PROTECTED
