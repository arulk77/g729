`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNVHJbgeVOieGatx5DeSTHU4Jp+4WzYIPbws8HjCwJ8v
h0vCh5LdCoPXF88PAnQnQI34bB6HVhKZ/KsikuMbma8U29Ufb6PH0aapMmwBeOlJ
XN18GKZiUl/oS7t2SIl0HeKW/6dJkbs7POFpVZeTAiGDBHYU1DB1Rpl81kJF4ypV
vAWl9zSc7PBUCLUQhDFZoxB5zDIHrqAXs5dAaoWRGFd+R+gGkH/0KQe8Wb1a7BGl
`protect END_PROTECTED
