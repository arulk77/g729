`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0z1NhbAKtbjKu8Ea2BO4ud67Db7sLx69VA6gXg2DhJojry4V8FK5DOgyREFkelzf
hzpnbSMJjPXCposMpCMFspfzZ+9+pb6w88Sz+NEigWLXVBYP2FatYFKJc5NHkvL6
vyJ0fdI2X0MIG818KU054O7yzhkWXBn3h18ilt8wnCbDxkX0fRYL/8JTa7HDM1Wy
oQNhZN4vk9eCFj5e+k3WUAsFDeXP1b0Wh3KJxFomOIuONI6QH55tsWdJ+k/L8wzY
rKggob98+L/2Msp2n1lGy/cjvnduVpDSIcpt5ekaKkomOXbCwjSUNNFaJOhaN6Va
yXGKLrOQMPe3g6VF7/ysEEeMMoXiMzR0mCIJdiKQhExIhDqFXTQZIgRKRLMkCrZu
Za6AbSQNmz1Vo9I9XxxT/F0lKroGaUiQFid1tcdUo7Sn65Y+sZpRkQ2E/1BQTKwi
WUBuZ3Ko+md10oE+LpmR20alWYIFPraMA748rX2jx3g=
`protect END_PROTECTED
