`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCtG3aCVvhDHVVXy3rJ67USJpVvAsfJYwqYokrGHqSA3
Y6V+3rzUsFMgidlQjiZICIoP5l9qhegECbZMXLQD9HKoIqDh6MldWfMhA/+8J+e+
oVqL9gVEZwFBhOejp1YzHuoDiO66Cm/5d13dh1PbNvi/xfk8FOgMDJnB/43U1HaA
lEK7kA8/aDEhlTyQ4vZD+g==
`protect END_PROTECTED
