`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKOoj04tVP5BXhImpOnld8NgzeoWdBIldjcU2c0I2fdC
EiOYqOfcBIOcLEx8h9Q2xkNO3KOGHwIpUOK6aji5/evt2WyN9aauoj4chVDxROxg
wVZ7DS53oePM6uQM8/gICE7NSIeft9lzljYI9Z35+jpmlYfM94dWrUErGiYi+6kz
dSozu+7khD2Trqrk3PcEe9p4uCfFPxLgf4rwDvysuePC9cagT3mDsUv0z4basVS6
`protect END_PROTECTED
