`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C63Ffc4VHlFJwu/zF6/OJli5IdkgntGa9LiqhEpwYPxY
U4t3MpSrOPjmHzIiqkyWZ4HVpelveLb7q00GMSTdr1a5xCTSOdIp9fyclM2h5fmG
7oMzyADaoWMspnf3UJaA1vQhFyaigDeyoDe5TWiHQL44txcbLH/h1FNQh2uuMxf2
6T09lqDWpdqjsKlkocmEk4bjnxRMeLwlHMdLJp1zrE4pTpnePlV2uMn+8FfXduSL
90DlBlvyrrcZHnVs7GH4V3m6r12tvoRiD9AE3VIxacsxGPpf7A07cDIfTmZRwjMZ
6nNg29WOfsPaMCEbL1h79XIkddu7F+T7NmWuzjII2T+zem8XUBOHvHZ+k6dMi2pv
NwP6C3gcnMrQ141yA9HkAk3lD3Sms6zes9dkVf+K3xojj40I7LuXB+cHSZFGz8rh
VHKfrAkNK9GGuC1WhEpHtwqHZ9kgf2GavYNbbF5tlVfdIPBchZvR7um5Gcvhh8a4
zFbanDcpERUvbtA5XHXUKSoTQBf8U2q8jRGEtzfyF3jIWgVE5lmKYFEgAnLs1Yha
H8X5DzLcrQxIHZVgiH0eu1axl18ZT0WLjSC61n0uwSthcJ7ABTDzYcYyMQTjcNdl
Z0O3TnglF0kP8nAFtr81LsEecfsWGgYAwWvWC8SrRE8cn55qJvTvCYMBLQU+dhkK
DTVmA89+A4KFztrnKaxWDP+q+9G94HXItO225rlorTSuLqirLsdRJIudAEOCFWtG
uXO2+5PqBVKvQBeiMlhb8lpN+OL/y17IEvSjm3kmzrj6f3zxxJv+pTvbN1RIAtfL
kr80keZs6TAW5JFYBXO0y0QWeiZ0H3A+1ShLHEoi/XpjNV9Ad5j/p14TSNroDfXn
t3DlGd2ICk5IHy0ey4NMFe50gdBxZ+4SgJfx9Zz5y6gnkqBSvPXN2TITEFZyMb8T
u1OSqxjSnp4DvpYcms1kIp/ACVIbJmHjoyEnJlNZm3K5/n/RPLomlbXSV8zFkgss
vDGsq1dKs1B5Y90A9rJdKWSzmkbwNgCODTAndPewno1B2PCXOMzogny9CEo7Z0B0
cHC8pQg0RtpMt3Gs87uyLzp4cpBJGPAbxy5Mc+zbgnUcgdPVdegiGpVaIXQacxbZ
JVfEvhBSTV5dJYpPRZPNIRiDA7sxsyU2ZvR4uToEODH2utu0x/vFTyXdmDQ4AURJ
dV8tSTZjCnJIt+AbDD1qnuVPdbDJvQ8eCVD5w2LjmYtbzXY7K7CzIs9o+f3N1fAr
GUbIsqjEqVPaAjbEjr50/5rXYRdbadfLeqElFGBSucqBwtgode8dzlKhFOIDQxyv
7uv6Wcsza7rWdYeMYeBODLzGFlNHRX9UA+WlM/OPEkFdPRCvzj1ws9bXEIfI0/8N
yBHHIotRd+yh/vJs4PRMawkk54HDsS2Pxbpua4eLs4WuZJ1QKnyxlShHI1mye7kB
hi3rvPWNMIVkbnQcdOc24S6o9XHxuGFpvS7nNt8vuHjBQs1/6gQDlzx/zilXyUeI
q2XmLPsEK+HxBNotbguieXMYGnfy56YoeYejb6XOrqBSbziVCbKi7nfG181QBKmV
8GrleXOFZRkzjBBNSe2QSWwvBOJIvJGj9boz6n3F1y7+zidUVe3htuF5oXy4r5kd
gWWjKcvSHI95cQiKzNThrstYM5zeOlw0+hyIEPTd2ckuTAAC4mYTZPLqGdtztsU0
aPG0M9C5hJnOQ0pN5cVcF3qN6PF1x8EeEEzx9IteF4ik07ZMmC6TZw3ciZMaIEPH
Ip/6IitdjFmzCs6b+u76Ajyt1RkWi4ZM3Xk4/bS4BSSuESeO2k6xFB814Lo4iwRi
BqojvW2jgobe++inkdqmv6Q40b12iZM61Ieze9Yexmorz2WAb/LE2YrwtqRiumAY
p0zKGHrdKtcojhDsPMzcX4TRpC3RZ1xgp9fYpqxewf4Gcka/mY89TVf2pe+Tf9xU
RL70119g/+CDnWsfYm5+1LuGMm1018rJQB6b5uFG+S4jvThZywAKaKteq0couyck
hzDdf+20B+sjT4BSa55hHfbytRlo3/XPAhe+3zXRguA/Q08dZy5X7RtXP193+1AJ
tOYe1gtzbyOzvmq9zGPW57yWSl/MADeyZcWaHbaXzjiw3w+x6kwcsM7qHbTKDTxw
OiCrq717gzdhWG196URLF8Z/gp2kwjuz8VLpoZY8BGhrtlYPHCZ3WRI9zl0rdO8v
tpIO8kgVaKB/ECYW7J5oZ3Dy3cP5YHbo6WDRJCAbUzjM0DQaFYzPvDghfLq/9Uzy
fQbaQinvjs5NvupVP3xaSTwjHyw7F0IlleZjEBGZkiquaGFOOGBgm58WDBVI2KS+
vbOHdbDJ2dge5jHAd+//PQaC4BWlW+5SceuSOCXzi1R/S9g9tmoMMIoG6sCl5mar
OdRWuiFqvm8vqmG6wZY7wA1m+LgKRxfVxK99+7X3bv3VH2zmuVMLUVAmsseAL7dg
Q2QHFSx/9H57IctGc0sQPqb0x60XrC54jghhpb6NFdPqRplFHcIyCgbOyL5IB0TL
KSJbnZKNFm53MmYkaXTw4fcyZmwZUpFWfYgVIE4vk31nWDhzWvpXBKgmDOJUvcYt
2w/TA/z52jPEbhfviQCjIutRniGejZUqXuJkH8w3+D2OeuVxkGT+RXWUEhtaLVN+
SzqA6PNLPwdvIcU/G3aNDqzcjaox6Mi1n9g83NiGiNrepDmoUf1033dPLwCbfPRy
AXcQjraZ364+IRIpoNlCHabbohlx7SqcDkcsVatqLX5kEgtVJPQ9QlWSBYPjDXx9
nkkoWyJFxp5QOOJsTBGqWFZk5NrFlk/o0BiCGmS+VBfE3Hv+jRdPCeGCuS4A83xA
CerP8l80tLqVCzmiQsVICXhMidzakty2BG+w81Ob/Qedkj4WcjC3mPBxT3kmbr8Q
Tgg9V6eJvITs+eBXjNvOO26zkNf2D8Se9YlyFtTvTctDkGG5muKuKikc8/iSxAZi
/OW2spK8pEBmYn2t8Id3SlDG7DQv+dx9E2DPlJB2Qbf5AVT6dE5agZjZiwxTaglg
VAtOgix+g4Z4+4wtpLSo3ELFhpsC23QNnCoiZeTo8QpY+w/MOFxTkwYNMUOSO4N+
4dASI4VZAKx5SQ3tiPBpDXhtdUJXM+wA/f+JXsMbaVYrOwUNTKUNu9mmX6Txu+LO
1bkpL3x8Fw7ipogTRw56kaGvbUaahS4ONWBbf7tjrtQzNkXUh0blq9ny+p6EWWmT
hNddJyDRggWByK6p86uIcHK3n3IIymq03882xYcEuOCysMtDtY4JZzuDGZ53HE22
vVD5hsBhdynfnbEmpTw7CIv2kmQe9IQLNG0sFxvRz54slcGKtggSHue2mqVlfwTe
jmhb0kD47r7P4BBrjg9QU1H/EUb4PSJw3UPBJkIeQPmXpMzimQSkAoqZ+sWBvtgp
Hulyx2T+yxDmcJUVtCSTEwg7RwRKysJouEcyzUan7osRHV40wkIhfBaeB03ba7dk
H1b/QqlFu2MF0KgVDF40wqKQjIDLFTCk8gjStwxdYdFIHlZ6KskVJVST7oNwh3oU
WhGI/vNq3lI9ojvIp2dB6uY0af4yLbRrJrD8BfAcin6OSPr8CJGBYywFP8NmQX05
fu+qr3+7Qy3whkJbhNtxo0JrAmm8uvDYDLZi6/S21SX+zx0cDY+P4NUV0LEBm5n5
76kBhkIPIcjY2oyUxrOMut3bXOvQKfCfaxczeq+CM59UUg2j0+/9xXqDJr0Qfy5d
Y5rgzWNOl8HRWgxxLRq9dD0ewyBr0Ezx8xm75IFgBNKr4Oc69jli9e/9cRxbasdj
cjaLeJRUAtl0ge1E5NAAuKvwaH4qjmwEB2yTwzKGQ9kpFm2o9Os3t3DhjYMjrHII
Hl1JtV6fCTjN0lJdGWJ8Azrr3dxDESgaqjVqJcBSCEvoGvjEI6wjuIALiqEfWbBs
rLQpl5IQANWY7lVn+n0a8qDrBWjgHL0ylkAlu3EZt/AJBf4pPYijGdJSdPOa378D
/ueQJZ9Qk/yh0kle1OD7OOaMBzfTSe8phisCqC0I94RYRMtdH1s5M2KSd15MYegs
y9BKMCwxN4LbVPnfOa+dgNGgJniiuEi4PUM+QSqW9Lmui9Y0ThE7ro4SsECS9G+y
UmCNkuEdUNhijqpzlMibTL8ZABwq5SOeoB850fuDIQGCl2WG0Ypux4UrSeHSv4X7
TYIheRu0az0WSr3DJPiSb2Gf/9NWW28KyY+mFM3m/uRr8Q0dsjdEp6c1CTILXGKY
ub1qgp9HfIRZAeGwKHIYtdgVTQd/xd/tJP3tEBBWkyMrVmZbA9VhNRvf38O8lUox
DGim22gI45aqu3K8G9KZPxMnghIng2wGo9/Lw3/snsY3Vg2jEyfaSIG1dekoq5Ci
pMYP3Qs/elgE1mltX09i3g26wTF77JnLm9XXs3+XYq2BCm46efxjuu7dDdBAyAaf
z192YMsWIpyu4t/+c5vCtNw17cjk20tlGP7FeaCzi4P0YHQRig05u7o2Bo38U16f
x8/3iSxqODUR/kjvNPKbC2r60Drc3E7s9aUVpX176F4J0V8EvdHgTbw8M8ZuSnYV
llIFeCTufs8FrH39qAKDqyGCOc9iSaddyQq9bk2gqnzDrcnrqEPkRHCl0/hfiZC2
dVZOs3kemhg0x14mTi+o0fVYInS6KXLcRwIgOtzPKbtU+yLsetfs3CN8Cqs+6KzB
4EeXkrF592NB1gZJmiDQb+HWwF9CmKgbUW+j54l8eRRE0xsHfDsWeO5RMrx6lS49
xI/Ipq2aZZDCfCCn42omHkNtxG9XSND0yvtrf5IlF3sHJps83fBkSlihOh6C8+6t
xaJ6VccrmX7cp4Mqn6uG6X/s44nQ3P+PFejPsQVz8SePhLKWTnUrQM41EQ9mqJdv
OQUrmCCum5ElvzpNtEqkvUgv/1x9Hb5KGpM+eTJVFj+kp5EMC1wITrR4iy8LDe/w
fdQLkHvJNgX3E4AC3vRhnZqTD+1c5RVAfUE+S0bb8VBuqVUuLQjBwiCMDGkG5f/w
tatzL//kQW9sldcMXtM7+FH8VjyYxayOcaS2tQT+1EZ+RuTD+V+aElJXKH+T+bLq
k95rj36X+MtbSNSN3YFULmlRMMFBoRyHjXVAVWP4pRQsVsHMQSXwSaE/mk+PuTKp
itROO5nLmuK6xm1iwAnx+JGnwTutKqY4Ki4Xr9PBY6vzZpR7LsNQqesRnze3qhJg
WTm8B49ldjv4MHEIWcGIrlp/XD0P5qMDUvFVOFs0gwxYMUH5+1feEEnVbTqo2Ouh
DfVGF6sGrRLiyWJ7WXdgkG7Zgym05x67FCgLzDzW458dFeqmaOC7hpFT7BzUojaE
d3VEblcWkWDQPvp01Yeq3HqUyHRxgQCXAXM+C5yNfY6jROjVtLbx41zBTPVCYn6v
Q1n4pNpfDUu1CgvB6Uew+ZuEhdh7c+gz21kCUz7CPPyljq3qvrRd36U85JBeOM77
6k1xD7bDyWWdtCsGn57r/SmZLjHB5Qt65ZG4FQ5biybEkDqGJF55fqBwkKY6lYEb
NDWVm5mNpWxtOLAdfSt1WQ==
`protect END_PROTECTED
