`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqnMi4iS2KckrFFOZBqFHVgnfPsEy7b89Yr17cBKkMHz/
7xHXDyLVahliBg5SIVY+UR5XTsjldDoLhnHDm0cEVEv/A2d7H98OF1Wgd6I3C8OG
QrQcYu/T47PIzKRmq1rT4DKu08JvTMryCAt78/avGm7U7x6//rjI0jObqWZzdZvo
/c/gyq4/quucRRdLRWG8GabsX8/2vQxkr2L7ItfDf8XJy0kCikByp2q6+j8ZN8Qf
KDpV1yenR1yshpU1Uw3eyHkZZvgRnTSJouUjKxv8osgIkeS7FSP14PJOKJKN7kpj
`protect END_PROTECTED
