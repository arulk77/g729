`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEFLt4fn4+QG5vBbM+f7EP79X6u0K9EH8tiyhpSPziBH
uwYSG4Y61dZkFYHnDQCi7Kr4V80duAwRr4NIKFEmHShZV3cBdAXp6hIzg2c9NODj
z1JpcxUfsV4dJiVeqoDjREjMNzmVw2wMHnk5Zz5T953WFRxlGYkN0lWocCidvykS
RfODxq+RtxEx/gYxXCOvPAYd9Y6iago7czB9kzJ/ytwdbwdpMptUnBqBpOtnyJID
UGQJ8qmxroKwlknzTrQoDUW78uVIFHCFdqOy2bL/xlCa2YV0y4V+t2YGyKN9+hbu
fc8lSX2iTIRzA7nvvLN+tg==
`protect END_PROTECTED
