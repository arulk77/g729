`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CXDo269tkFVLssJhCUcbkcgIbcGWyjVb2ysgEX0OqcNpovM6Jk+063UCkWvgxO3I
zraT9z1/vAmvoG1QCTNU2NG82EBQQUZ8XdmxgKiBObzKCBQQdhuQt1VwmQLvpy0h
F+AWnADg6pKc+eaHrUiWUBLKIuCZl2kw6apaY4KMbJqjiclkwkhnWs9oMpQSekwV
`protect END_PROTECTED
