`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ccdR5dVryThlu8DItRO1UyeRwLZ8NnWDUbZHRsbpkUWV+b6Po6qgqcn3M+GGMNTN
WljDZh0PjSR/xPXlZjqB1TlrNU8ZBnnJcF7JsrDxb2KwBMed4olHwz9ZDTNMDCE7
aUVhPPwU72FX1V+rFDzSzvlQXrPN6DtLmevSNR1ESmyGOpG63BPWUJu7R1fKzemo
yDbwMMP/JniQdn9EOWY/aox9DQi+QVbd3K90voYWk2ioDURVSPnRbMR1yzWE4dxS
bd+c+K4pqJ3Y0Y7u0DyvKlPw94vs/gnsflR5RMqZBgQE8TwDfahjbWJdrZR4v/3n
rKxxftXgt8UW4Dsok8ViSTB7NdotHLs50I5nUXU+aw4MmQnXHmUlqTqAl8zmoB0M
84Eu2CKOkmzjqHrfPkCvU3K6Wo0JPksGiXYpktnAeXmR/RkbLS21BW4Nqf09/uxz
4cgZrUdYbkn0UijzPLH53rhDP9iRntBCw9sjBGU8PcwkYQ5+DBXvLAAPD/uLNL1N
r4jnEOp/sPR05B0Ni6fOZhfQAKJYqqhDaQt2MP5rOlLCU4d4815ukruEvg+Hz3lO
/My0kCb0j728L5S5KIxEDHhBwUEjla6vqD/bb2XpnOgZ4K6HFdMt1v8rAiZJQdVE
S7/MtpqFWh/oytuYJVCIZw2Ky/WMQftrCskoiqsp/gRywerloccctRPk2DELX3wH
jBNuxdIoVk/ILdVx738EoVIWKhKJS/MNntBVNoOMpo6DwUiJ1ApgsYWm6mNacu3l
siOjlFzx1zNiQm0Fx/VisUDnkhVxB2DxXObyDxre15pWL9r6e4Uqcwj8DUrr1e1c
yxRgfILKJBUl0HL0RQnaO+CfdjpL13JH/zZ44Uv4P3g=
`protect END_PROTECTED
