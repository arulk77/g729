`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIp4fZIA1udqaQjQMYl630CpIk7ccZ9vk8r+0vyd+QJv
RkMGRgcTHl1sAKfuO2Ts/7ByBtAJxLR7pwvEPdIY8maRgWxs/VcgJhLXxwKqTzID
7rVEo/qqVp1ZIuoMjfX8O6ZPYdTv882l99bHvIrt/gXb6F85y7oeVL35Td/FvaGB
hEuQaO2eGW1RZyA5C5VIQmFEbQLDOoVnIcZkXyXoypvEacB2pprF3cNH0pU4g89g
PRVmbStcygr3G5HGqn+E5ChBfrcBlQAdTt61Y+mja7UNYYlQ2Y4a4RPNn8XmKvgT
rsu49bOsH+QNjGyLB6S2Vg==
`protect END_PROTECTED
