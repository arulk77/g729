`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBTEVH+A+VIbZ0UtC4nPtho/S4Jk4xmuKOEGVBRJDIG5
37VKellvxJIe//+aXb1IDdTAi66jI+DE/4i6amLuDdjL64xPl3f503GZHLiMUUpW
2qbWfsP2r9OV+Z3YouTeKA5KdiArYHDlQmonV+zo7u5pOBLqeQKdsRQOLayxTFDO
ZfYbEzWmb/eCDb/yL5nfRRG3ra2erzeAKXaSHSy3i+U=
`protect END_PROTECTED
