`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9GW49965FO5VgHOU/lIe/aJ5cUEbycwRluGLdlbWsX+S
V8B76exeXnROZCYRhuOyCuNXbmzlPXrsQ6ugJBXPIWGk+NrxSpNEyvmfbtdtvfDB
m8fne6/1ubmdOzhd5mSMccatqn9Kbl/hVWy8ygRhKEIENNyD4PgVgBHvj9P6Zl+S
q6NwRfezut9Nc891bSp3p5kua7LYTbIyOlb1we30g5taMOQuRU7Nei/DFIuElwF7
Gx0l2wOZj9zkmg4uyxBBQIkOSKIy1QGb9EvxHFeXJp/HNugDIrdb0V6WfKf86sxn
TUQ8SyJUA3SsBbfJ9aggt37DYM+tavzl9dOGefdvy0AXNXkKUKcvyzJwCuAh9LcS
/ktkr9bHvO01pTJ/VPl0MKLUSlRuJuPxZkz0vJoQpR1I0+MN4Bkhbl+Aa44QhYhv
aKXz9RiLgmaY91WdWMZK4vgnFKlG8NlDIgfPcXsNqw3sXxP0R5ejeo0IKC0Lao1v
GJylBK2U48LJKFb8BhjFPcm4pfPiSsIhqDDEm2naQ2LdJ4aoPH0BhQAdkCAc328O
XLvujPCh61hNjFGJXFltr+ZtTkrN1zOfF4bCrfDiriDcMJ06mqdhWagoHuYUFL0d
ESDKMkvZAo6ea1O4AxhYJu5f8TaqyaT7DsoWvdGSqJHiy7Cc3heCMNBdRW57L7iO
cEc1d6yz3Ul6CDxtt+YuwIcuAA28rcQ25FP+RhgFlml7MEMyJetyJYE4KdpzVk79
QDcfBbGbjCybnYqT+lA+ZS2GnIizM+YIwp/rneltIfXk2q5JuKpHkoPCdryABvwk
Cvd0U2mUIMvceqQYJIHr7ujLdyLfqimmzNMCRPhVkUdLC4diKga1NfebTsFT7McV
ZSxx6a5QlZVXf60EucsO4LXejUsKKXI5ULs0qu2CHtSRrkMWAInZ7l8mLiHe82gl
qK3741cSaAp6WM2is1FkZLJeub8CAshzrV+Ewx8cmFLBBvCzjOh3mO6uV8A9R6fz
DjfTC3QRSaCbm8+FkXEwUmpVJxEp0baMe3cZ6CkvFkXTzGNZ3WqYzaywjRik78aC
Rp39KGL+WxgI7dfDb7BPmPe/sL+LF5ujmLBfWqr0a+atNYx72lEgCveJkiOPW8xK
t/N0hGVsn67H/GF6YfIxx9OTRnN4XH4G847zFWQsizrAgBwRSb1+87NN3UwBtieP
Bukez+BEjwKzVClWxMjnL37V4Y4yBnauDAR5PqlBgGIxFDKa+5vTjyXOOqkmIsv/
Jh0SkjY8FyPE2boJrqDVRp8pVjeWIljeKkb6aMGPAovDXGzw0wKMsu+RG4mJuy79
JwgK2HWUVHgM+CwXyryl7JwHJhndv2McPAd1sHZDoR074iPliwqgCgyZda7riEZ1
WPcVNvhR2Bq3hA6W34L9GvEjH+HtTXYZKJ3Cf7I7/XM15Jo7HGCJNwTWO8qtCiZ9
Kvozp0VK0naNxERQxmaVis8KXYyDLKQq7RCE2ykAe48FygvMaP4jhuw7NCQBVZif
WYJkPFZ+K2vqq3OEuv69Foo4A1zXRy80Qr5dofHfAypJgaEQPbIVWoB9JJWlRTOy
zI6zw+NIHgFVQnhTf2uEVxcm58itE3cHl48oQir14oAAEGm3mgnpCfs4RGIa1Snb
VYfLg6SfumlV4NtoRWeZt/AzsRie1Zr0YJCyfQF7w8ul2taQm9ejiFlgsrkXAh4k
2i3y2jhHG6mRcDrSKfUvaooQ74RP4avpLc+sTStbVVaQfo+iz2S/UbfgBv7E449w
MY5Popv+twiAHvO40UDrUXnWVSNzO4Yk4UUwv+djQb456/jvA/XpLJUIz1VLw/qO
IUgXrvlanHQ3ZDhrxwMse3Aq1l2X49DmN1EYYWSrS/GDl7oEZOTQel07yrOAA9es
RUqm+wF8Db7qFIkj0bbv2eLU/tOGjvP1jF9C4audMLpVzCaEPwW2EGrsU5BwCIHC
dalEbjNgWHY0ZbHL0YiG4wIkvfxx9IupWghsoEfket7Xzn0xkP6xZSEhcApjTQyc
hU+A66QFsz53tXDwueVNkYRJawqWsZzxOeuJS8PHnCWD9Z578RLxa1OM3j0lstH0
MzrQ4CvZSpWX0rqUCA0v66wJxjZnew3oLpsvS03YKubbtDyAhpYiCLm3NrXWfdHX
21nTNf/MbtuX2Twxy7TfutOKPuDNEJ3+/ha5dIBLr03vrOcM4Rw6JtbeEKDKfU46
3XUOlBxgvN6Su49UgF3CMchHtS7tbY/jkdUb+f1HBnX+L81d5abAM0kCsO+qIAM2
sGo+Cxyx/88OV6r9Q3KgApqHKzFKUVJ1kTEAp1V6cscnkfGEu00ZQ6KEMIKMpRhl
UnmHnaPcT5I2uLEBYAklR+oOpcG0KkNVoGmp2mfH72Xf4ROelRB5JRHhbxppUNNj
7eyh/hXIm0h8hzuSRNx/IsWIEfsA4GCfCs9UiAfqCzMZey+7Mi7fB+lUs/BoRMld
JV6taXiXpcSqIdTVoqHLKlW0xhWB09IdWs6nqSEfuUuQYctEyCFP3s4RbZ09oZa4
8MVeAoWBN8Y9iz4EGMObeQxZc3hUCywff0+Xi1kzRdZ1tFo+mrfquN6bI4d3WWXf
5o1UfHjC3yY90ak+ishBJRvJhgfHn6oPqLpox5Gr+V8i+7DFfdSbGT+Yl1ylBE10
2mkIpdE3Nt0ux/uQOVw268NFPNbYfKDtthZ1iInncCP7mNi0lCAqps9PfKT39nJk
dql22GL+eva3rX7ZDd2dHH54Qi+XvewwzXgRPCODNsSDLi+4wsXzsyWSqHHQqG8q
zJ8TPLVpGYwS46H9BIjeHI7SwDE+eOCuvCBwTjWF2pZ7W+YcJgstwO8KeOPDWzE+
QdIbOwvTRgIXiIVxla6QXz1Qefd3hFGcnEKhlxHHnLgwZpHEHnKUw0CdDqS5pjFM
4W0NWNo/mRzsEaDk4nVah4oQ79UZtVui9RxkJsRML1Pqato1f32EqXUyzMhlsFyJ
PWP+JVWaG5EyWaGjSnZ2d3pjPt1z5Bh/9koSealEyWedNqopC3gZnTHUnvsgDJxO
x/Fd4d56qT/37L/kSbGsiEXv5g6pvphI3wcWkAo4MLnl+OtWwoTIbzoI+Mlvq8eh
UZtAaWvH4KLrmG3UlSKvKlTDrR+HqVuFkLJKt5yAUF/8OBhheqnXc7XYemBuN7oY
CYtVkCaTbHMe6tKoIeoyUr2hiiiBA1v7P5SAWiZWY6/3ij49L24XCB6f3kE1rLcA
FZYqGAdQxEXQyXOrvNFN+OgGB07c+vTPJQR13VHgJcE8RvHTVEhatxytkrpPiXPn
nbJZVfq+lex027HtWI4XvLOiB1aV4DNGbKYN/T0jBcCxneKxQENRZxqPaxE9NgAS
xKhCnIQK1DyyLkMOrUK4H7hZjEDBSYxvQUnyqc0OSz5A97Si9FfbE0LDMOjtiSYk
/Grnpuqa+FhSp+yWUfI7Dhd/5YOUF/3GaCbmuiPjopOxNw13I9ZaygWlsId9wj7I
XtgRAkw3Ili/mcGgGkLlOoxOq0N1QpEeTFCGbcaARp2B2D3JFgoxZcNPHYYM+cIs
V7oAlV1XrJDpVeF0cn5SLUZrK+ugpD6dCzUqMwW4oZ4ip2luv0vuBzFoexnalWDO
N4OTBcjzx9Ln7kHE04rRNEVJ/4lhUrqVYu0/deAEmsFc33306laP7VMXKhjjHfHw
EUdQYicTOskGghTk0pGpt7Fe0Nk1p0LVxu5R3KhVkN8HqeV5KXu83LdBIJPmHqDX
QwtlGOhMSbvwxDsgMHTyeUS7w+XN7vBN8sjDTwCXh5+GxhddRg7SlHGTCNXd9rB3
cp3Zdk3/m+q5zUQSIBnEmZezpdoa2si21LlWv/RYR1LFh3M75jSpoa7StY//LC0R
xz0EcjJOVxxWrTMM7aDrxiQROM8smBIVA7oq8/fEtvVJyE3CR5uM+y5fTp02aSX3
ddMRDsMEis3ckkuR+KEcmYUqnvzLWZPfyzlgamG+UuYmM+3317nfnotBnsJWEyer
WtQNIXQ8StsEfNKFzj7uA5A8aZq+qCJbbN/7PKTxJkXB5zHHYmQQR2Hj+NOBRRGC
JrLRjdYV/uTl54bNQKwewgxK5SLha1kpKl+ytZP/OypQLswZ4AjdHpIDbIwjqOwK
QGIX2ovvduBliQ4TtBR1iEwTM4drytq06UoSUwRjdfgmjU4lwjNgk1Fc/oDPeTrs
H7HybijyWufkJdl+hmk/XvEl8t474w3rCz1gvw+sYLBDsUfQzs07IkWxjLV3iUQJ
oBaUc9MAoWH8GqCwIxqVxcYSK+c54qmwi4QPp5VQ2cZOB+ri351tYiwQXriCnK36
vOqgFVPvKSXIEClvmdUhdWtBGOtD4sXM2/sBerbRL0U7LLzjlGatKDIsoavecRh3
G4PrnFEjgoRhSOXZ5NeDDwABk6+THDayRZiPBK4/gkafu9bSzbUoHT7t+VcifBER
g/fDnWmx7itYeQiRcme/8yeQymalwOuZHpl4LlbXZ6VIrd1xGGpcU+PplbyHvU3w
czXeSpScpccyu+wzZLBsJ9h62J4zZWM4d0MAc8BkYXO44+kkMTaAHeGLyzxaNk4/
HllEs7rqzGfVUWKR1Ln75u5UdLgmwM1EO1k0RMRIoEbZVYfmxNWwz1kVVhWrrycw
AjE5i2r++yD6evX/BgyBObbdzNkOx6pxQ1eOm1XUfCftRpAbE2D2XTnXhx7GrzE2
0EHK0YV46ACR6iQwwsbLolK/2iOjr+atSjXCMtSrmZsNa+2X3RcETraSSr/AjT8y
aHx5Hf8Ep08mGphi8FH8m8Fe8fzwdikDrYbv4717hBna976UFelrI2XSnNK6rgN5
l0+MQw3FFLTBTHCF6JBb368Tkhn+i8I3bqIMx9qkFI5qqkBDZ3/+U2fmrxZj/RBJ
CIsbEg0Dc4MeKfxl7eVu2+LRSN48a0zBf+RcZAQwbdhXDMN2556LfrOOgmtomSvx
E15RwToYjDRx6gNxzUA65pUmUQZkTQiLAra853TT5DVkl8+GLjU5uXghz+6bwLBf
O2N8NluvzYInNbNgQJYbVm3+BfzB9OPbCj7WvNmqDWrehcVOpkNORsf8xD5GCf9w
9faOQJIGzPpxiSwIldU2K1eDAqBZhIqTp4SIhb69Gml3OuaYKzGQzUFMCkLmoqnF
Fk18apJ+BiElSjy+UqmRX28hJ0YEAmBGkwXZJSn9arJFrqr3y3JgtTMi2UKpJ2p3
4Tiw2UftHNaKnLJJ+j5hjcW8S9GcgBhsUmeHn4R7/DIUTqRoB5cXBCokG6xJ/qsD
fn7xvpLuxqB4FsYV6cM8pFxMxG5FS9ewOsIAY3n84lLInrZ3zmUig3fJmkLE4eBt
al8eqOGEBnpFaqM+QeALMDdwcsHO8juAi/2dsDaLzfaVDSGn8xOn/FsWIeesHEB+
9ed3/WXXmhUIchEF52g39yKP10F01qD6srIN24Uodrc/2NjplvGNzGtCHo6FU7Uy
yc8fC2rRDa2HqHqdSsXxlgisG55jCZy5huh5GgxG7y2TCv5+Zsf2wkjJs0FamjjJ
BO4pY+k+WmjFx2koita0DvcGaTZgIkN6IjjysYe7MmfZHEnLy3vdRkYS09j3l/fD
u3KYgfwfbHZWhUMcx/5N13R+bD0oaJIjtGGYp6Ny+HwIB9FsEqz4EEAHDDVtN1wK
s4fM1QzB1AWC6lJTMDN/OEnvSAdkDWN6bOPX2IPPTpVijAKr3mZpua2h+3BnDhBe
Xq4aaxZ6liRbAft51RFLl/Bo5VwmZAQbtfHuNXudRB7oxWygGUtVk8pCFvx56/p7
bhRmBmCniBVAoqAKlqOVHhW0tSJKAfK+AAw7UG7owsfd8CX/HN/xxWMA+PkYKfGi
zfDjzfcFXD5Cal1NN4enxEdzelKBH7unYUsaR/kl/GKc8l/6xIYknTW9uEkRtddC
8jgeO9N360NMMxCUhL040D7Twu5m/kJprmyD2YnLilnAbJLs1w8b1D5UsLVSCWMg
b/r39XWzcg7ouCGu0DC/3Ql4DKT45kaHtZ+3auGhtmHqwz53XbbFoa0MkIWKQfNa
EucYGISKVfpXbvFSq3z1Z+BsaCx2koZbatpyfsVKPVaEr3Ggn6guQLZpjfgUL/Xu
J/zuA/b7RYpgYGhWoqZMY4hd54E6/2n28mhV4knlGdCBWgEktlPuIAsTfqmIQHt5
mMM9A61jCcROJN3+5X8juYs5bKvkzfp7g+knKbtvywxniA44nIleJJCSCyP4YWNd
9iCdUn04Tay88T/hfu4JgAJj4/s9YKbu1KJyOamLifcWtt2/AVrBvMJaxcaPNfTY
ylAOKq8voTXo+4Yowx/+EA3yU8/Zlh7w7qsvEk5bRlkCJ6hgckENMGuVl5ir+XZv
19jMhOclLLixf9jYpZBJw04dX9ELrWGIFT6AFn/r/04TE8DJ5dYoTzcLV8PxUHae
wiLFrvfL7JwexQIw32d8X8z0N/Oym26gpjbJwp2kEmDHqxiLyRI1DAcX34dIdau5
zN5jWeESeUWyE4c2igzp38dX1TUirw6LO1kzM8yovNut9PDm45W4YqSfoSjCS6h7
2v2J5jgAVQwoTXmYKMyLRORI24ekKiTGbdEoMYvzo/L25Zj45d/o1GFp+eEu4eG7
`protect END_PROTECTED
