`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IpKK6ZJFL25IARZEAqf/LHiGbfy/CFGwtPhiBGnq/u8I4Cuh51dRLwDpCjI5zwi8
CUSzQAtdAVjz4lnCX5/Kdz5pvYT/+4gnRfFJF7oa80wclS9mrB2/xTtWyNJbG1MZ
emek+AlTZS/PINppj8j24Yqol4p6L3Ff5Govd9FWieB2NG0VsvQEws4saHeXKmxJ
`protect END_PROTECTED
