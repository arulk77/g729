`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abgHLOtHdiU/NB+8CqDdXZChYL+Ivqh0PqJPsM22m+q+
La0zaOiojPYsntvo14w+YdSbPx4NKMJmn3JRSltHiiG/UWZqedGDLOLonkEtpq8X
siG+f88T/MA//Ao1RdIF8CmlOoFnPW0MFiQsCbQml3La7HnhYx2GHE7EcORoU6S4
r4JHqcZTsTD38PiYPxzwgI377Bv0UHP61bQzhEoWa7c4OQKhiGGZBsAsDovUS8LV
gxhB7gTAzmwHcXPwfkWuBBVF7HJtrlQM8WTU9oC7P0sbKqA/TON0BDADiGc+3D1n
J1fmII9T73d9K39t4ZKM0sBfGSCgtEkw/JSY9fmzuVpA27xVVSHO/dJP5a/1nZ/X
ddnGb8H8/T08MWflCf9Bfv3cP/6p9GasJmMhZTOFORYFOaTY/Hcdvg2cck20MUNs
v2oP1gEbtdvZoXAskhVWAQ==
`protect END_PROTECTED
