`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xALrF484BYPn7rpxIrTAAHhv9psg88j4bxFfo3qg3a5
ALhUnzQTO4CQDXT3Vj+5gNI8xMizoHI0XQWWXnaW/040UTjPWAXiDKwGW78JmQc4
klWjI3IZTMvM6ZPVlT3D68hQUM7A4itzNVJZexHiv3EAyE/897LbktqzHjR2ETpt
NSTTmKpGFuferwB2ZULC8sby6WJN8gsDQr3mwKKPHoneO8hIOemzDfrltgE4pd48
jeQy9ut//0ia1yezpLOKZy37xO6+Fhx598NZ34vn1yzJbgxCUGiqkbYuEeweTYYs
bqQqolIBw5VMSKh0LQ7zlXYSDHY6mKNJURgm5s+vNjVaIcbpkpEpNdpO1zE4rAmu
qThPu1ERxs3t9Iiv2QoHUw==
`protect END_PROTECTED
