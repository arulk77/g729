`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL3g3WDTN1iS/rnfepiWwqOrQrPYawIfTNp88v7Izxrk
fiI9zxZwPHlNnwrEyvGX5PzkZdPvVoGeUX0KiDRa5ecNqkzuR++bfgQF3PgVXK6Z
FdYLHajSLXyNpjEcBCXZzuAkNdfr+BrxUreu1KF3hKcwXE1XyML7Ea0twIh4OUET
SYppvQB5nHi3Yu1E+5T2muLKoIn8x/xNEFH7+Y1jZFDyBZs28cJfv4gb7eWwRn3e
+MNfAfw+YNjP664P3LZfNkAOXen5JoD/S52Ail6zBHflbWZ1flnZVGjYcypx2ile
iTOG+76jf/FCxvkrN0I+zLT+wpW6P931UmrbQ427B4jldvjD8ObbYKL7x3Hn7lGP
cNYYBoyUviFB0EAawpm8qNXEg6aYRk1DUP1JHmngJf6PAXZJOS2zCTsShKYXzbB+
xJTNrB3ji8da2FEVd728dvGZAWnr2BPbKwffFEqmTQhH8tAw7HUrtEIQx66FWW8V
hNxRDVJ4mTgNuhm1MEzhh3e/Vs6k8p5hA5EtNlla3meuFiQ/W2GeWiQCHkI5Y2zt
`protect END_PROTECTED
