`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxJNWo1TdrNtunt9wBtLZ7ULVVSE8UQSiKJxIZKgqrNu
i8LI84DJNBAcDueOMudY0jVOXgFjCF5oQUS7po44ZGjduVztYcjKcVknDe7sfnwb
h85Xm0kbLvCVN11LYhVvGpFnVHYmEaKI6wvkUeUDQT9OnpZ93KzE2W249qhfqteH
XVxEghdUOK9I8w0MYRNfJML/ez4Z/pJmklRgeBdv0H5cs73E7DcSXqWma3lntGGK
nPRr7mnlSz1NcXHlv9pN+mnmVfM/kCE6FLoaPFwP7F4yDvdMwSrjagWJWLkqzQwx
1O5YiJZ+CFayd3Etf50Q0W2/sMLjyfuYtMiFnAgWw+1X8KbCRkxglrwiyzgtthuX
9CQImpSpN59HVhdrY02yThJkdXwt+3Tc9AJ4RQdh/5XQbrgaT5bdrXbQpGqIUkR6
C7nJL1S7MA+MQG5fxcmlVY6UMu8Zqc64cGFTZ13fTaA8J4jW8eipleWlxV9R5tA+
9dTlIjCAgiMofWyNva5gcGi4CBcR/XhE8426VV4qpf2ZcnGsSYMfeFFl8Ya7x5yG
j5hWD9r729Ox0OpVDaDS4zE7WiSF5EH7bdmeunRQ7mdZKdiABW8AmkRNs5pzAWld
OQ/ZpKNT23L3BSV5dOWC+RSOwtWhSCemfc6xbf/ennsS0ijcsauyNfncj6FOHO+s
hlN0KH/uuOZ61fll3Oc2eRe+U17SXfZyqdqVGPa1mwJ+O87beSxygGjhoBtcLIn+
nrIFMKKZQJcdrajHhBeQvVhnHoVZEAs9zSQRD+YRYO6AHnx3tKzwS4sEO/Zmyolo
vVnq1jECbamdKksfLHBs9+SzCKsyxZXBKWxr8aZ+tyd/7WYxL5ID4Wf8X6VYNSl1
cz80eLoUZt0trIOU57qOin/vYTaPTHmkULcaDl1UQNvbwrfVFc9ex8gVR7Ai2gIG
ANoKYIQKuVVlffjuy/Nb0huLjkViCD2R0iAgwPkAJ8HnHKiYC7Lf33xlCQri8Mdi
ZTC0KFJypmCoy3gsM9m8lbduGHR09pzBoYNZzUYTV1cQNaBLkOzKTYjQ56EM7vUQ
OKojHCZISM78qfpOCtKJzTYrrnAUHN27gk5FaFUyp35gDlyM8C6Z492vvh5pN9pe
MXNnuPLEQmM/ocH+J5G3a0hDDiOQ1ktotJviCrV9rEf9X99uP7+CFiJBwPLEuLMF
7jrlgceh1WVDHxhUXDYjSOcDk1Ihzj4N1p7CSPlMWaUXaoxVwtabuSZd8SJmeKHh
/MzLW9UsxDPUMMzAwYf6T8SfE3dRnZqUxRKwrLZAxLyFga1rB0M4817vX1NYhHD9
jlszy5Ip+Srbr/y2DitMLprfSPAgLKf0+g2liAv03OxaG2Bto0oa3xhuOairq7Sq
AxA5U/TJ5ZymMEGl6h2F3tQN9N+PdbadULARvJGakPVYZGZsn+pwKj6nRBKdr7Iq
qZ7Z7p5tzeWsSKFN1/A6xqy2pRtZLfKMDbtewc2nsX3CLKOCwr7fr4zI8F6T3hL6
5eHsIcTGxTSNxDMhx92O2hEfbh5luJOTohm18sDQPpxDPluQu4qc+h6+6+Sq7NwH
uvIfsWmzhd3vihLGr37to/KCwWgJbUSw0TIWrfGZs9AyLTEziCXFK3lei8u+23VC
y6HraL1BEB2lQQqlaAiClsTsNcwYzi1h7leW566hpzgwqzDPpJwIY3m/z1so3NXo
nfr1edTVoLAKvdSSTEiuiEulvrRfoyuMgqcarcEXLJV30aEHf1HiYTHhTODE0PwT
OozDK7Bvsqgn+0IpEbR2wrhI22HBML6xsoaByaKz3/VDwqbJUFNcHNyZ5n9wKllF
YQWL1rxNW5Gcgay0GtXWTlNlbNIxqHrxSp/pBuykRrE7f77hDLXoZPQZWUVEBUVF
WfBQ1eft850gBAnU6YVuAi3YNsEiZEFXUNVygORjQzQirTlC6E91SgPITPVcOP9I
qazz4hZJBePi3vN0d39EoQLnUthBnutASqlTOJlEpymagyThJf2lF02w0atsLB2J
GASV8Ub0Hwvg6krn2y6ZPksNapqIejHV64oXXNVUjlVgg2LTu33Qd/deJM7NnCIG
Rml/QKAWZaUpjgQpeJGaejGq/lBRg8vKLxTxg27GmgQgJu5buAzoOsPf07Ov3u8R
v7ij1HPIaQVoxEBEB++YDiIqRCF4u13wjTEit67tBLXWZLOPcICgds2Q8s3omK3C
CbQK3DdJp9DWgGrcnzna4Fe2vDfICY0lWpro94E580V/IgKuG4DQHYu1yI+LL5A4
zmwhAwzTskpQg5JTgVpAodzYKP/S5Emho9HN1wG8j8O7l76pbC6ZlAekSNGiBMUJ
OwFhpy8JsCSDaIOOJvtAP1xAqXP14bFouSEy8+W9UAzCpxS5lV8FUU+1J/lUrSDl
IaNzOcbrISTuC90mN2Esxue5sBLTNIxqmxxZJEujaZZhprRV3AOxPREu1lhVv1YU
rMLO9z0xp4QWhTr+KqzVi13TzFyeSoYnGpVqgAIiI9KRIbYG+TzxJCHVDLVq01gf
L4PYq78EymN4p1Ki+rz7Fvdz1qXVBxNjgI4SwPc0zbeGHw4QJjgQGAsHBMaOLeaP
i3GDduYaPf9HXWDUY6RtzKzMSN/yXDjHowTU+z7kb4E=
`protect END_PROTECTED
