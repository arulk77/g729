`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFeQvcAfPc7MqbEfADNqfSX52HWwx/rtVaIk9lnuBiJR
Ge4Mq3bQ8d2/qEZ4UVN/8Iqdqw46Qkaj1ALzgrgJQpzZNPoh+iUv/k/W7rZocRs9
LB4dcHy2eIJYSAE74bAgi0reKiKr5T12JTflu7QH3WXjfPy5ZQ+LQHWZoClwwJPu
DFO357QaTGiNDOzfOXHtAESGQC97GdWzFlrr/GJVh3m2qqEO7NlVbPDOzhhonZ1N
znRgzujsz9v0HxWw5F7l8+g5sbESW2L47UIwiReiKmBiCnRod9iQPqfZJhdMDBMK
14WfFOT/qG53aOViL41DDdWsgwii5Jp3zSUbQ9abcuGl1vKCinuxZI3fLvcwAAHV
jsDcEFfDjKCiQjdWKjXBjEDuatr5sIsrxMfW/5STyLglFll+KEC4AtH10Yet1qfe
WUTjse+KxSGsPIQWm81iRBufeGhC7SA/OLic2iUmzCQTT3u5BtUZUV/+Bzxe+0h1
DKfZbuCrqnVd2Kzf9omWZ7+oe9ffcFJg8UEUwbG3sh3cZ8W+jDkkoSHnmNb9c/zJ
US0l3g6pY9x6QIvABr1W85uQY40MbzKMeqIDcx0ckfPs4ZkIQ0Otpx4PTz/7ZdRm
VkbhEzKmUntQMn3xPoY5ukMseBWCh+BZqitMVRNhBg646l8g5MnawAJkcRvvQCyO
t+rGKKh4CcIpXhD/T1yipUqSIBkhHLHfbBfeyvdQ7IqYnciKVBumARaJauTi7vXg
lAgiym0rJMs21fPnUYP/qC+V7Mk9HKjHZd+9lbGp1+6EcfmGUU0VVglRDawcT6fd
CiLg8HYuYnowzJaNf9OmQ9UK4Q2sYm49eD2orqvIDWlg9ySpmdQ9y+Yjc659/aAH
5MMK9pDKYeP0t32MkOW4TwNGhGKdD4s9PApiD5VZChU=
`protect END_PROTECTED
