`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42cYkd9Y7pes4gOqODK2Hji2s9LqsBAlGtCrFTbpgtlU
7DaW2Sn1k/SJwdEqpKd206DGPT2dLI445jeNQfe4hEGVBQ2O3d8N6GezrZ5lc8m5
BWHSjJYxkCuMzaSkcqDXbiLYjHFA1WFr/fy8zRvcZsSmrha10dEdruTk6iLZHCBt
KAS1Yiy/U7HCb7XdYCTDtUoyy+1d7JExH1SSRPzwCYfTPCrbyiEaCqQ0Y4NLAYBL
228+9tj4HZeifdnqwYcpw/HreX/iKyGFgcsBYxtD122J2czO+82lLDnFBEtoYO6q
q2KKgwAjEi8a/LC49qMScg==
`protect END_PROTECTED
