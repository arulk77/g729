`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLzUNA0ZEVpL+247LPf4vIXwHQH/iClPhPFZpKMIbarV
Np4p6DOYi+1/o2hUjPwmMllHjkyx3lqNT1hPtb6iwSMzhPQ+4nWfNa44ycEhs43p
kQb48jpeEV26OZ1A6V9DMsF5rWdTV3/RtyOgvS7UpVF277EvBmjyB7PEr7TAndpA
wF8M0/4NLc+s2WbvIdx9qJQyNisytB1aLzm6WDVt62p6H60+kYYbBMy6cJ+bvdWG
Z1Ci18760SO6S/Re71DxNECf4usDDe/sMEUIe0y1WXXdTsYpPWK8fSUEQgHgDkuH
6HK0cBMBPE08W1BxxcaxFQ==
`protect END_PROTECTED
