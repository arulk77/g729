`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
m9HWH8CcT+nKBernmW/uNu0r/RnvQFZC80Q1oIGiQKiqaSe6P6hTAjUwn2AOF+04
wtLzT8IUFVBPIEAV4TvngcqsWzF/lkEjMhsx38TMezVomwpWnCn1VYahOevCBS96
kCtDwnQRFVEVFa9GkuvsdZpTW5G56gx3rHWMroni1lzVKQMLNHqwBkW1vmIGEamN
KlWRmJTtMhTXwEbKrtm0rMit+TqyxeM+LZI+uiUkMBgUFnme9NxwSYeDMGa1UwPi
64rNfytp1Wwi8iYsV5TidORwYCt450ge6YQyeQOwpZpeAzVul4HH7ebPDyxDDx2t
P6t4Y3uKuio7U29Dg6vh+uppPeGv0r9tJaJNleH4Nnk=
`protect END_PROTECTED
