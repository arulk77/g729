`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
F/ZPZps5D7MCvtpKef1G0MQ+qyt/rWI8oOvLI8cxQ0k6vxhkxN/G8flciCYA5LvX
9NhNJkzS33f9fHOXcjH5qWFaPhdsgD4LGceR72TwLtzq833nk2WyVc71VkktBid6
Ot0iEkMmppRL1iC20+Wh19Us+l1fV/Q1VWTk75B5bWNODuNB0/vnktwQ+WB5tE2k
A5BTtJ2pNHfDlQTyKcmrDSCEWGsz7W4PGw4B/5hk0tPyFIAis2k4AdCAJeyb+V1z
lIHsK/jKcsBdT0sQV4YMEiBMcMx7YhcdH3sfcNIwEYU=
`protect END_PROTECTED
