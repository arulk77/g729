`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1afGrl4ddUYi4a/t5ofS5FtUFeWwSQAn3sCTvT7p2wf4e
JqHe4AlMBbbpg9Abti8ZurnAgDhdDlJWEaPt4jrldscbbG1bBlYNeyUhhHvs3hwr
YDkoTnjeOHdOcIW0wJ5qQPHgvjfyca2p1o582WmTHR1Hi770/BDK7fr8gMDZ+fT/
tYhcD0LjN74vFrPUwFNIbDYE7Jou0Tj03lClhKrSxlRM0knVd7aydsbudfycsfMT
30ZNXosuqPUvrj5bC6MWvoD9z11mY7hrSvPG9epCvaXUg/q7HrMnyh1meeTTOBnf
kV5cWf3/UvVZdyPdWubvYBzYk2mbhDtqJ6qCSYhweAU26ve5ejvYKjYOVh82Kl6I
5ZvaLITf1+/xoW3oRIxvhNwEA0YLQAm3qdlMXv3ibGeJl+ZYJo3Fl+9YzY/9IiM0
qMD2Pf5D4WNegjybj+AP6C7zSnGBvwteLxV16/m2pVFbMa615+BgofyAP07mvmGM
FUjlMRBiXfN+jpLbNbqEvxuRryRI4n5SKWcWrLJk30W696IcUslLaotaVmHunWjG
VwGFGBjWUD2X1phL5io7d3nZji9nBdLUIDH/KQy5B5P7qJJDHi7EVMkUtQ4L3BJf
OddfymmlxWYynWyXDrAVFwRbZAzxX3nju/Qkr/5tcOUYPK99QLo3OqaYosAM8Hbz
NbCQ5VAGwyuB/db3ioQHcbCwWw8+AhqiQX+wL1EzBrjn/EbDXTzQo/dGoZ+YI4iI
IPrg/CkOWl47R1u9kE3yhRgp6MFE3hwZ87DnnouSyfUbDJL8wIL8ZAEzhV+Z1iJj
LwadZygSGR8i/1rFrzzrrOdptJfItMfpkaTweEhFWsqYHFzWr3fhFH3fypNBo7Il
yOrSPS9HSCih62wk8Ww9w2xr9SrBUXdsakoJMdFJhH1qSUWDSUGG3Vyf+xEOxhUy
xSM0Z6NEBfcJxZ+Eo4hROAGC4/mlVQ5sOHd0+OzmCwIK8wJVz3PIAqlJsiUwQoAs
ce8tYQzT4qplx2biQEDvwzw335pigwEgHsmM4/SPkRYxfp8SGDlYrAQuYvohI3R6
0Il4ehRLk2P5vtUoC1pKTp+bqNQ+47QCNSllloO5NrLZOEzIfKd9aF8tVNffs5Nu
SZDwLyO1EQGXF5+2ccouZv7Ax64Pbo/3+zpUlmJl4PJchlyPnWdTKy4KvV8X9dCm
AmQwvwaeM6VbjCm/e9E45brOhrw4oktHDJaOWx67HsA2rjy/8QXUcBOnOUtuWtNR
JBOqw/x23GTAda5uX30vzvrgkfDFT7FJk/m/plO138xj4U6yPOBpB+XIXdhgFaRK
TDs/lBUIK0eRJZl2ILIiQEaw/leg4EzWgtJzF5ZwuVqi4+jy02PsurG6O2TniU5O
Vm6muxEXnx0eMsOk532IYl4S4Z5jKshBBvUjk/Xv3LSUNtX4kYQk2cBp8YxIEpJ4
JxB7T92Zvv5jjNQ8rzBAQk9HSjbOg/Vx6kPpxcTqxCJrrNOsB5U3Az9OJ8ABlioT
6HeRp1VTYJAMK2C1nxuiqUneh9ZLxluzV9UDR8wWR44cMs2gryuue10FPiYi/pjv
rAcX+AWtoY22ly1cZsMBrPZiqsLYII3nTTjGB5HbVBWxVp3KVMw0EB7sj+4XjqdK
Kg71aQ4NHgDWwMIQNukRJXk1aWFZZ13XyuwCyFvqZOihQT/MILk2GFXS1CZfIU1m
JMo5gpw6uVp1NAm5HAO4rp+ROe5Cea7yVRh26VV5kTtKOj1JnBrjE2zCDvWQfTQL
ioW+QnnMZ+hMyi2HrmD83x4OAvok++6y6q4payByEC6Mvb18LEoGmal3M/iMn1di
jOC+R56TBN5jj9h0Eqt5lfccSAFx+zhL4hseSl9TOThqjut+tv7gHo7WHJpMMi6g
Pfk5u15y++sN7RYhcYZcXb/8EE+in36rbG313tiSeifMCWBYXK/Lm4sghhvxhXFL
21UWiL8aGfs1aau+BQve8BCrVZEw3nQk8405ltSbpYc4kz1Ylq6ggyN2mwyymLMk
BkdIQnSsC1B0N29CjayVKQTjhj2KeHCO5x48h3grFHO/ORymciO2vrgMdBHS5exy
e/nsFq3AX02RIQ90I83Ejii1jvmWPIM4bngQz5dwLuHyPHAG+is7MSTXOIeAxdKM
WlUiRVRfAOfnuNp32MLHFL9RzwYJyI8lJfNj+m5xp4lstN2qlNm2xXisSbKmb+Xz
N9MQT+PZgm/mIFC01LdZsge5ytHwI84W+Ydq9XKqa9p/cdek8jvSn/TNjkLadsJ6
ll5XrrnjYJnk3WwvgPW2y2ysvES97TjJTOAXovtGDRdG7Ov9Wo9EAXCG4kJxzExW
ZzDq+LnYB7/NG91AyFYlS5c2KQ14PoakDtUPpxrIhQEcs9+9s+YiUiIaFB8rgz6D
RjXsUXeg5QwxHI9GYzC+M0pmswJVb/Vb0TXpMiVHVOeJCM4MG1YpsABRKqzdwfHB
iqz6SI+wntZZqq71D+Ah8jWCKKGbU3yGHTQs6eizz4D7X9tj+fufx6ctCcpMGABT
AecIR8yuakKjTSPfMM8hjiKDHO67mZ9ZU1Z9mVPlTR36sOKkE5WEr0XY1YXDc3FP
Ko4cvYstb8ZX/B4iKpRxGTjuhLopysn0COB2/f4bKwEm7jtfW+cYqSybf2h/sFMp
+fNKewwsr7zgkYSPgGDjSpdFSv1O/Hieb1LKvcPvnvIbGByGxDfBEW06e8HLPehz
O9tvzb6ejhxcn8hpew3mWk2Opnn2KI3Yh1kGmx/MPAPq06+2q/6sv9fDIL488wcT
MRfwdjBxoP96jNDHjZRPxQ==
`protect END_PROTECTED
