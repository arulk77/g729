`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+55FHMVRclcky4KNcvUwgOGHf3x1DkPJkGbkQeqRzgt+YbQNSFncHUlORJCV42SJ
8NbZ6CEl+hAW9SlziyReKe9WVP1eJfLo8ADxS71i/GVBFQUyIWRdxlFi4iNeYdWo
ZRV5UsDlJbIIvlHwpwGOaqucF3uv7FgROKvH0NmqR6IKHN4LeSX+8glzIX37zHki
zV3yMGg2czbP9v+Vts5xqIawb9dMNDGTZQQ8okSWtW/s3BUgN1mQDzwvKko3fMnX
lUeS8sfHkHf5Y60YcPtXC2gTNkVxW9pZR/4t9QBTxxWkmi+HHvGxI3GWTamNl+f6
bHHh6ZiMzg47stiSxJrTt/PJY7j8MofRt7KkavBXC/sU08v6ZLIYmV8Yqx4Mf3GG
0VSGCVjpfrK1eI0iZnNSeMtKVFaPnB/Bhg4QPiHV5ps=
`protect END_PROTECTED
