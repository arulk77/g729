`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePSbOqFX7uOBkF+gEMRx5M4yWr8GFC/kicc0pCzC1vth
7qCr/XJb1JbXUOR3qeQvOBWRZeAgnKC0W5vSRXjkvejhCNRApHA8U+ZSEmsLa4bB
YqLLJsX7mZqY8h0LXWXwi32R/7iGgy9drjAILd6Qjmz0Va+qFR6ZTnsNaoA4e/fx
TxRgdcg7HCUwMOxg5r/QF/d+Sj7+7+ooR7VD1XXVGoiGwp7FGVfupIUbUIrjjcVU
wZFVwnYduw5n8xvcHqXD39DOWEKgvC7GzDR17QERHxIn76RHJmLwNRUh8wwS7PlR
cgSZqdSk+A7ak1tJWPJaOYhnNRut9/BqutzExtF59LYn9v1WZiDF7VMOLSxkP4lL
s8aOYcxcFgtRpjy57Xld6iXg+0UheFHRyEApqfWZBhZhxNy0QsiLoCairr2tdMQ8
0900DlMiPdTUuuc1bPMSPYZYzyWuiUyUYYi9yQ7D5EXPivubW7eQREwcX1nFhHn9
xXix5CWHPPIbFHN9mQO/AhZZfYhyO1ZrD2FRgKcszcwkRjg4hwqHknyVg+rz7rZH
PREf7rBqf74EHv68hgnsxQ==
`protect END_PROTECTED
