`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK/slDY/fRQtInPziDo+6uKb4rRVXZxRxWxwCHTlvVwg
cCt5yiRI8z/3gBzjYOHsfqnTEgS9Ztgz10aNstgRZj1FXWuNbiWUo70mLjGIs7pl
Hy7WUbPlxFzphqTe8Xs4mxOR8XJllqHrq5J2igEsjow1AOqjlXDjRyOrbYsPgOO8
XEUsrwtlWdYXrULW8SBooFQSbAg456Lnvya/XH1PaXtkA603psvVAqneDBE1Gub2
6La3uqLWTpgD88ko0Ncefh6Hb+u/AmQdNeBhE+66+AGwkutsLJzrJKbuLVNo26lX
liHvu+uIRo4Jvro9ykUQR11/jMrJLzzbUfUT51dYPWcnIDTV2hZX/QjmG304KOSN
`protect END_PROTECTED
