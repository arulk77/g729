`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN4qB5INmuIjDynwWam1HvgpEvTxJyiLZa0TA043/ErYf
QsbCH8Q17ShFulmhHJovdf4c9GDSObhztNUC18pnRUoseCPb+1U0Hxqw+KsmDPKE
79D11ple3o78/JpPzm/23YDFgMj2Tnhbcl896bGBXkPpcjYPHxnH3doIZ5/iwGEn
8HaaKeHXcXTa24aiUq585cSxuop/FG4aZVRY4k6N5NmAceyU60Fo5esLrD1kfn7t
mw7EAjaBYh6o22h0XW0nHnSZ27f4IFm199OwHp+NuPs+sRWmWNlbNlif0VP5VsuU
syYHhh0I8Vm0kecYIIz6akeyEHN/3A3N5ShNdBRX28C4AYGhA2Oyse/s9lMhenur
`protect END_PROTECTED
