`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI+dVY3SC5HxpbCKn/LdMgHZRwmeLgBQG+S+oMC15nTe
qxN6iPRlFdhE6BzIk7wX2HA0PvvrhBXWl/B+hx7KAmMgfl731eTI1V1OAMPj6aJs
ZUtH8+JuTx1F11uNs2FKJoz58Ye5pxeKhfhSx4t37ixkjDY+muPPHwGzz/XTi8BL
GNsjmiAw6dyY24h58R0gvmVuP3AfLX3TcfmjeylC1iYSZlhFIJACKFdCQ/AxGNeT
yS7o9HYGRAtd7N1hTEcVQunOUPWuWN7p8HZdDlBYrBOjBj7Z6yL5jdUS7F0s1XAM
7QuP1CsEYuKDnetbBDTLHNwyCmcsJOQmkW/msL4BX7aQLcPVTgv115l1UuZIg2JN
WRSyU1d+q+IXIJrpi/SBuwie8v03wtSSm8Mkg39hfcCcBw2yf1wU2wdlj2Lif9oi
WC0xVyNFU/XZKd8UFISfKF0AEyYC/HMspbYx6cX3yMuBNoQf7qdqCh06kD8nHAtN
hasEnM7IZrukVP3Vxo7WNoaed/hArabEUYyI3IeLq/5RfOJUxwd/zdtzl2kTAoOC
`protect END_PROTECTED
