`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hVeay00deS+HlrmTiEEc6PL2W/IS2Gy3+kdSBuPR/iplJqHlrbphv7XQCyD4X+0R
nvUT0SNiXoppTJZS9e04+7XuCijI6M6ihl2LgDkI1bBCYqXDX/qm97haNldfoO3/
A1suc/OAjy+c76w4zuDVdkodD5BIBhFc1HO5EMOl9lqsR5KKmWCcEvxYuZSDBd7Z
97yYd+7ZvrmOHMjkIyhEcM7AbVKx+FU6/XZ2EgrTqur5DPb5iVHJUF7mSJ1tvQ21
wPDl2hfSHfV4BlTKVEbKcIJoQ6SZF7J+mcqEqY+DCAi6IpzwLLRXKc5OxjvVG1Pq
mBL2879cFR+9GbSBmpu1EQD8H4BAJB6XsFex0ROHpufb4Im78v1rerwd3ArzJANs
Iq1meFsNSDi+QrW6ARRnADuNBc3fs9f262cFCtnV4+I=
`protect END_PROTECTED
