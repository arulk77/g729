`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yQYn/Zp+nG+Ap0Wm3ONsBwDvQYVgc9hZpom4u8nBTte
QKjyTWiPx3tGvlSvGdLh39xp100qkzzp3xYYm8pBkJ7gjAc2/qAgiHau8D2ZhF0t
FPMht3YmXMsKaotNPwEtWJDNC0tZDyIQyhVkuBRqzzhhbub7w+EzIRURY/BwQA+C
wdfzfPtwNotplzN3lnYVhxZrgZuT3HQOFml1+TP87iFA88bblBIKl4knNd+83Dgm
EBTl8OegL7wzTI7k6ZZpPoC3HFZv6sl2zm+76DcVXUendBrIrX89bi2Jilaoo2BL
rWxNTUFfK3T7KBbJIfU+V9FLco1hVVDFf6rL4IG6cmvgHyJlDu1yz1I75w0ly4vl
zWT5wCU0M5irEBrFkTa+yqNWVyS8XXRkdC05DAVfDaSRQNxLK4DUMFWvNX76t99i
7ZIEbXjyr+0zqxcfRqzXOOi+6nAixuYAb6xJd0/j0LpIMf9uLJcnP8tFSqhBMUaG
`protect END_PROTECTED
