`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C24dD8Q9AIaimXM+1x91Nf19lh/hGX/9Qz49Ju80zFVW
tS/UCdnbAC+iiM11huxnwvfi0dta9IeEU35+CQMaNXFCxKGyn3yEHXil57FSg5eO
8fG5DvARxFNh17Rxq+Jx6gcTWMaBwzp3ZToFvvtr+/oGLSw+GHI5bWYCibQywdHz
1GBperaf/q4e63DV+BzQwKfp/BrZpXBXBCiBMQIoohe7OguY8FgF4WFJPmD2PAT2
/yxvG/Qme/OSW4LIY9oa43fCbANZjz9eik4zRn9t4/QrkEmc/gcAbjlxVPIHQsc6
wzGwlrG5g0YErJoyAr2QuIrIhyu7RaQyXn1rK1KJ4U/21eOWldmB4Ds5sw1yppuw
qS6x1WdiEOLYLn+TMrIhK96dbIkh3oI/mGPgEIWtWMmHxezuj1tAzjm37+gWYLhQ
6fFPLB4G0Wqeb5VAPJ3hzzNBTpq0otDGBPN5nx1SQxWHIJcYRQ8Yio82XGyIGEGb
tuDMB6eJYVk5bCBRD+YKF9BXzLQQj9FohHLsYTsOhifAd6ifL/bC1Km8a1T17O3U
9cmdqf4pLDZO+xUid8LxCPC9U28YUXTlymxZoL+CT1hcD2Q9dffJuiipPSVk26ig
uLHao8FKHrB4g0oEE4CEwn63I7WdasQ121wQzu6s6LQ/TsIK/8/QozrBDHUf558l
XOWgC6+lQxkEeXV5r3Lw29Z1JqLCTLQf4/vkcrgM4DyIMv2ORm5G2tIvQZw4LHpW
anTEfM+jqDz1VjZxZIRELmUkw2qbe2Mp9Vt7cLZ4Y6F8OkHe+/niMLks5TV7A+2F
nDopzk8YrrB3iejQTNzAxVxyN/U3/ZdPeT/gLFUWGCsjgWA3p1b5r5ZdCIYW2KWH
B65gGVziEIuNmX9UzhIHo8CI3fD+GNa6B3y9TVLZMbECr0XHn2O+euYhzPkaWFYa
mIOeApwcYgxwCFmzGeOXuV+38DE6zl1TT0yVtU9Kq2MS4mZBHtaFtpYasQ64SqzA
hakwJ6YCTnUCnOL5BGASGFmovnihmrzo03gpQ846Egeks4obi+TdEYJCA4r21sg3
I5RQY6TMljq9N2G8qsXzap03yQ7WPom5YrA2Fh+b7y8vrsrASrsGe04x5s3gFTB6
LxOKbgDqDJ2prDXa/5SF36Dv8br33nGSvT/DhSb92DVwqjJukBMgl1KxUhynZdK7
AzlKS8CEcOkF4DtObKPsqnFhKTKbLetifqHUJU1Dh6VLF7RinTTfYu0DNrecHQMd
QQkIJX6RIDQ9LLh2HBCYVJiX/oWeO6pQ1GKamcl5fSq3uinRMc+L+Gnfy0rxnmKW
YWTcSjFAmR+ASF9y/epeLivuuziMTzlKMoryC0maUCJw/D7WBkWhqzbA13InAPo3
vYXDi5cX7XGBR1fnbfhPldP1CsEW3L9AvReiLZdSVWXkRFa8ypnhzEG87fvIwnEH
lzvg4HELANX9gZyFFvT4ghNmIFism523kMOa6v3TeYEV1goqNAZM6TlfgDa+EiC/
ElnfVN1KKYivlrh57wh8vauQ1oGRKWQ8lUsD16G7VSB439W4jkwqlSv2szTXUTe/
7qmXXQtEIYvqBb3tayvgyA9g2hroFecAoOaiUXrNrYIsnzjKrvWVuhX/M1YZMX23
ITMzVjBL8Gv4lMttNPdFqcWuWuaMlD+kQqKRVzcjRaHxcwWrZyeMQW1HgHR092Ba
aSbk8IR9QNLeUCoBydEmZxwJb1cljHfoYadGfJLiprE6MTy6cUvxl5v/gyrN1kQT
GMCL8yLolMwGALKYpN4h2ICjR2kaAkltwVkq3/cmqxjMTdjqTwcEEIMYjEgPyUvz
iklkQivQdB2sXHZPnEcyYAw61tLtFL0H7s1kFX9bL/mzfspgHv4IzB5p9v1q8RQD
aDgQBci/Ey+vwDGc/COTX7Cu7hle6+YwRSY/tmB9+t3SVZiJNAhnHb5w4oxLDu8w
Euo4vqxNFdcnXyXw75P1cPth/fzFDEL1dshsm0cKfWBRVPgqdklJs+/6SPLKj/pZ
XhwzZFck4UfFwrLkAM3Hy51vYC/bTgCMBPla0wvzvWEe7yLfmw+D6Clm+BtQykYf
FWJnknfbiYtZRYnMC4/8mITmg9wVck1Ik+TuxcfzEZMyMCKnJMsfPwQij2H0S7PJ
aeDWcqW1n/icrTR0ACifmczJjyBJFQ/3DPOdltwtN/1bGHBItU/IwchvtdcAdnBA
pvphzgR6BAcQvu7NiDUvD07+xKa2tcM8cYlu3Bv2wipMgUqdSL53W/2WErxBXZ3x
flFAliGVnhMn/hcL0qHC9Bojg8oO97xUoORYm/Vd9MF8SKQfZfkhGBIAgij0+DON
RanBPukG/o3jwrunhPP9tL6zb3bQZrCyi7S5Qasa5hKMCpG9s2ysIx7z6tDFDLMa
U6k1uG1l0WVo+8n9INRh7nWgZtotouxgH8RRXABGN38JScs8le4W58xj6mgf9q9j
lPBb1UoWDzC4H4YSuOKPvqMfpEVhxxEgoWYEfjb16hhrQdlf4LwTSXkPuID1Si6l
BQBVBhpmMrg4NFmo4JvpwFol8oZ/sO9vOad958plcw/pcq8gQ82xzp3rhhQ5Te+l
8yD9PKN0dExBLjZSwHj1nq2vcy3X9V13LWQljWAsHyqzuGvYwQTJi9HkaZMl5UAs
+thD4D34iYsCid16rRTlGMna+04T0YDBll7ugjvG0DKhLwT6WsiHP6vFYsrQ2naC
BmydtTN/oN0rFNKX4D415GfqBhsQADMyw+r8FSpsKMTL4yWxb3tf/8uUVD/DGyXv
yJVbJsw80LHGruXJFWCdBx0ZFj76U7CPSI+RozIV30ngNcuU2V6UwSv1jETvVklJ
23O96qZJfNhWpyrwzUTsLY9i432d0H0WIDqF/ousLDyz+GuDvJbcijNR3mwhP/5x
GQLILQ0Uog7kIqLgKE3AJEavpEjJy9S8mvwuww0+SRKv+J34UPDbB43Ajrl5wnfE
UXuhbmPMssMjfIujU2jy26sD+RDa2s5CFlr3bNdJVELcu8UGr6JOVJKUAEeAJ8i5
+LVEyyC9KON55C5HIWisSy3+Skek6xPqRM6jPMsylmn4GPjZGyuwsC7UNBkH5qpL
s7tYwbQEYqRruJPoOb96dKULasjeFjwnX204mvnTHddu+geTHg8jbleCdPlBfEL0
lV8aLPYuj3PwsrNL933N0WTY2/ZonCOPr0gdM1jgUqr5WZIs8BgyZb3JJXvwp5DO
Fx1foC8l7J5yFmw4IDO/mnbUZAsd23G+63dqBAXfIcNGYqB337hAl3SPXnnhgn32
Mx1WXXb20aw8S3a+rjUAeSnA0ZxmxUAM1kWfywDV+Von2kMiykfRCbYaBIv/F4Tg
E0SDMH31YR7Jb0oDhiDB4RMfX88DZmpND3Sj1fDO50dL7MtgwhBvNSLwBRzhdpzT
rWe9wnZsQXNQmic77xcsbbZXEZFNjrxo0yIYuIbKmKclOKtf4p3uVAgD3eM++GMp
IjrCmJDUkiN+Pp/ktaqxkLCW8+l/QcJ3PTdSxEne1aoMNSbzDSdNEmN7YXgn8Qqa
yIefzcxYZ2jjr2Hz9t5mM7BhvfG+8Q+JAfZFGM/uR+rHmRZO6+FzNqROCW3TcmQD
JlV36ezjZKzREpJoFUh2flwOnZwgEDi1Xl+CNSJPqHNY1RYWJafP+dAj1NXnQXhj
F9i66aG7AFZfHlumFx557g4KMf7QNUTKgE8Fd9tMen0rf6r/pMfbwo7uFrxhD74V
wkH1piSDd1bauEupDbYS+SC1GHdDL3kP3LpFGGMQdGfIOBu1Pfl8YWMEM1meQLEu
WM8ZGROzGSTp1M5b7JcbmiNbewVuqNkRnLXEBxyWuvX0ODyk81LZuFTIR0ACBArC
CNAUQAKysnAF2H/wX0rWeyEmdCn0wj0Fm+u7n57NXM6Z2Gdko0HAC2PhKsXrGUqs
UAm2VFr3DYKZOZwxB27vzJJjiZLoJY3e+21mEPKc7hnGULDmVIRZ6GhPE/0eNQsC
r+XdCyRA99v9VW/GOM8eWeM+gYQXlCvbJuBo3+5nm5bblmYvd0b09QnUrUKC/QtJ
o4RpROVWgKOlEdZB7GGGJNmdP63slJO5L/CXWgUvp4uqssJ/1m0oPqFWUZn0W7ic
VYj2xKKbSOmibXmd7dbVdIjAB8XBk5V3d7sXIJ/Vv6c=
`protect END_PROTECTED
