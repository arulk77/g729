`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFFrr+Tvys62u9meqfaty/YkgWscuFxZp9Jvkl+Ld4/i
JvpP5xb8G+IuftzvJAWKDsdbEJAE9cH/4thJh3pI6sQQ4qG3teoQ+s61BB/+ysPg
nVcfGZGz6BmKIV+i70Kro5YmhX011SN2X1KXS1J2LZ0uil9VEF9hE+d0g/h4e82W
/8vQQO7g1ZBSfm5yXFxABufJTq6eKAP+2QoAuFqxbEEB5kesqiP36Gfz8pBxX63U
Rynz69CfBdU23+BJW8euZA==
`protect END_PROTECTED
