`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RjsvO2G1cMpQnm758KOobIYiSensmhJt9hDW+VSkvOVJJOOvBbYik6wNm9QWun15
i6v3jhzvrehWpx4UrLhfN7sKYm1qZ0WGciuvt5kYNHi3efeFN8F8ov64VMntyuJZ
uIXUKYrt0OTYr3LEdrJSDkBuZw407th3EaqDhuTyf6Nf9f2FKcfMOUj5MGblHRgz
9gkxP6+AuSMBB2YIFRgNcM3IquxVEOtz+mU/f4GfFvY+lXMk9za9w8LCLsssJWNY
H93JlmsYXORtXgJ8Eh5gVI377uOyNDLBZvi4A6IAo3ptrqYiYwNOGFYO9rEfLygL
kUKt/mOJAcdQsIGW6vQKWvfQCvP3bAVlYURY3rZ7Cuk=
`protect END_PROTECTED
