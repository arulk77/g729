`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48wPAQhaE8TfAeE4TmA06Q9+AWWO8wHfQu/Qu6xdaftO
Q1AEOo5FCQLS0oiUAKSaGQxA/sK/wfotm84RCqAoWk9H/zn5tAT0JixikqQSDJi7
sJrR1x+wurxct+zaBQ68Hmk7fi7tZmqyfwjP38hYtsYsm+uCcg4d8CZp0Wn8RElR
zMRtfEDHmUd42HU7Mm8ad4yWDx1QtFULCP2unys84gjHNEZikN+bINwmj9aDt5o3
8XpEh4f3VqFLaX3bn8SekAVyP3//0pNOpz069kLU/m+pmslJzOk1vrdVWFFVZqf0
7vMO5bre6dRK5r1a1pN6mW22RK+phm3E3rOW3wwMDXcVJ5JWvzOViendcAU50IVX
jqWKi1Em0WsdDxfQm80PQ9oNwX5dkoJfH2AjCa2RRhSeLW9hih/18oF5Wg03BMVD
VMa5WrhGdCg9LnjmvZAx6Ljw+HLHJqoHf2vpYiq7CAD6eEdkd+a2Q9N1jD56oF6B
`protect END_PROTECTED
