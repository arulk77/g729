`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZ3IX0GKyg34KCNQou/4/DenaAFuhaLTo8UBReSdtRQg
6IRQ5ni9knKj4V9SRLe94wfix6jo3BGR9kNqgIIxRcCdo+bVy310dQHklXLubK5l
JuwtLbf9FK4od8x4tDWzL1p6nReXAbnkJtWznx3ZOY1XJ7NuHV6CMsg4T01AdJGs
9BvbuPXk0miNmPZhelowNBlBV2j4O5NwzXWCDeblp2S9Kk+5AHNkISMlPfFjp2un
AmB2pyCP/M2xR+E8kb5NN1wXptqEBYtcSdHkQgKV1jVJlVIOBQaGJRGSmp7+zaBV
/eo4G3XJrLxOAj4dXCMKqjYiexbHS5JCPaOevyyBNzg5CRnCybVhWpdvxtRcYrt7
jWB8qQmJ3z7GqM/TO5sKqzridU0ez9cKqIU2985mI0sHBecirZ2mxM10HE/7Ft72
AY7N9tEzOxGBWzlQPKR6zjFJWdepL1cm2r1i13PoS4tUEFu3KJ6rYgAyhYtB+ko2
g4deUBdsnWcGphIaSNkP6ht8Qx331SUSF6W8cRt+o19NGJ1+Z6fEKgVYsoXwRIsy
LNtEcfyaHwW4Cm59AOKDCKVIVR1Wt97lzqh7UWkWtvRry5uTbCvtCN5L/SMseTF7
xizVk0i6OgkV+Icttm1w+EtRBzGW/swq+Uo8VcJcjzt9JaRRwxuS7ILVbbd5dSxx
qiFg7QI40qMcNGdu48vt0nabqddVuILdGfdL7bI390inHa5AW4S2GKVxaudXk+0o
Aqb6LaMZV3mTNST3TWKZP/Y0BCZP7Zt/sOWqc72r8OJB0YgMyu0wPOW+T2lzxRT8
4qom+XqMPoBR81E1dDpu5gEgKULgxIzC6PUsBcLshYDIBnZNeJioilko742AsFN9
jgo74Y/jZVzf8KSwACg/YHrdJR9Nv79S73z91YxIWXC3ZMH8SCt5ko1aAYcUPrwQ
Gpf8E+8COIURe/GCRrMa9KK6kCjVHKC++sTXh2ot4zH9lvvPTApgBFe3IOgeKdoK
uUGBkSgoatUAZ7JcziBussEiu9wh67HSf/v14gaX8MoNa+hv9xBL8q3R9UIGIpgr
xsA+pmRuVvQ/lbn1ZdmsNw50CqHQ/0BvOfMLWow9qLq+yBAG+nuqW6rXOxXgb6mc
jHuedMVWpvL2sXXHos+Rv2E0Ihlc46tCzsM9RWy4CD496qoUTQ4uw8Lp5AnXn3/d
TIureVeijuww3tnSBV20A5EtBPQVwF2hJQW5T7ijJ2Y=
`protect END_PROTECTED
