`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IlLXi50zCRWLJSeBxSzrKt0M4vQ0YqG4t3G9hxZ+5nQ2CTmeCYaK0Egrva6BdLyI
mNQFmk8MkRSlpEG6y1uLaq++6sROiwgXy0VOCK0yS18SBAR0xXyb0Qv189/96QGm
3u8ah7odZ/dWXRAz8hrujjVqa58tXUsSW4NYpCEsMMEqcNXXB5DK9Rh6WfkxPLik
fwGtdAXPO+z7PdBHqy66fBJLgWtIUOluJzfYhK+QY/Vdxz+D/a7CW0uuqRjsDFlA
Y3Sks0xFfzNdCbyo8MmmTmaTUYle8xhPFBwPvzsV5Zk=
`protect END_PROTECTED
