`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGj99WCdadS+yywOolVm6Oi1w41hlcWOXeSsnKk2Hs7u
Ef5vjCTh8ece9vhdk7tvknhdL1YtCb3BggJv2mnd43Uft12q+aXFHFj78LofT01T
hcFmquziKCwsOAekywOOe6M8lA0orKJ9Yhvg26cS25wv/70/ZUtjQpdgNmMnzzuP
LGRYYfOCdxhJJumRzBPCXZ33u2tF87L5HFurARSA9oC2eiVnIqFT5Z+AEm3jpR5i
ud9zCSwln27us0KL+fsBeiY8BUeNLnYhsjjaYkqA0Xn0iLO8kHnZ5eJkq5RA8rtg
5V5CZL6ArPCCEIiljVpcrJ6XoUrC0TizjfLrkm6PMTQwUhlYRKRNVDmowJDGwje8
fF0eqrwdKV6R/7+L2rsOHuW5X628hrIgCATBXlArNBCpq7CEdjyUdRUGAtiazReQ
UgjeEKg2JZFoW1kzYVi5rooHd/viXuBWErxDGmP+MCs3zd+LUtNDU5Fgxorx+eC+
mu6Hkxm8lD8YUq0DHnk/YD0HLqfUklacjXj7SNNHrmcuj+kq4nGEbCpAQyAljaf8
bq8rsqgsgzxm3JaAeVvTIGNiWhf/EMJi4HyStWfxTDxwLsrGgBNjuczWMP7WlPy3
fKD8HbgYRupe3nMeaNxn5leOezOyRRfgLOfV18I+x5TJQ2JKqoAtRm9xUYkUuu8K
AQvl3UsBaQ9D20ZS7pO1dxJMrDX16KkpU0CpaHmREUmTRneB9lxpin7QpJVOKl4/
HC1QlyJzc0io0xYQdXXruU1PRY67FrCVeV1idqN/A99o8D/0U3j6nfliYyc556HL
pFVE9xy45Ww9HPrjbSjY56Jzf/l76VfSn7nd/6B9k8kfPF20evfUciDbCxgtdAeD
KiMZwTjRNw4MBvUFnR3gaPmhiDO+9zOPTBynwnnAsGffZWQ8hBuAZ2Be6cKNRqiG
IUL7sxJ07xX5DICGpwgGbq7DU38cUi+01bnll1ej5U2LgwD4j/vwrYDr8m0Z/jvW
i/C6MV4D42tSVASssWV/r+NhL4j5Ybl5fDfdsdiwYPbjDh4nfjjpYS5YMsmvn3mM
fRm5Pnd03b0dTmTaDfjkmgVciJn6QCSsO8aCFo8ClzXCO6wUsyY22Q4QAt4TXzA1
fe32+Bu+eaSy/otc5U/RPIeeVExfRTjOYVxKqHnt51sIv/88rDVCMYdyd48IOY8i
wZWcc2vXNMDY2V+xH9WoDGokwqbj2G2y5znOXtbprGF8FXm3TvfYOQESJcwWH+hU
`protect END_PROTECTED
