`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7hmGnoyvNPDVft4cxclYXM8E5UdXfu4I2CzbPtmrfbS4
2qeJ68RunJsILBqazxVxrgsVb0N5VhoWNcDxAQttH8FUTK5Zj7GLfXr8SXfLFIAY
u515OR+GfepLyvncMIoaMsc1VhmhinIhyoC6gG6yHZFvUXCiXBls2fNLglRR+F+w
prnyDnIyJz/voA7QuLe13IndHTtE7P16wumRtVSOYLzEknNKCFjSVXl/r+QL304l
HGlhsTRzijeqc+s5ZtefPHWbc3xpd4V0eqtFNZzJNdUTgsOQ61B68P27cDhPHPJw
roDCWKD5B/mAgZ7vE78CaQ4Ux49wCiJNbT4lkqT5LeesrTIBnwM6eKmhzxCXQit6
`protect END_PROTECTED
