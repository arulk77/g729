`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIVbnp8hPATgxLKIvf9VQ+8kkLgGD06lwE3k+cbjcL3c
eGDev93NMEDiwnD87oRHvhwCt7mnoFzzVUbxSirGmt9DajYx9aq/DbGuGfw92xmD
vSY+Q3vXgG4cbNEwTSkNDX6MXHzKUm4thqbtR+9LzHkaPLb5+1VaIP4eqlXdAshV
LUBVnvsGeBuWb8UfnUncTh/kMNWAf/6WVNirzYRgnL5W/AH5O4QcztmbI2p9RSb0
98wdqJeaIUDUBx1v6d3lGEJecL+rmZ00N2PuDv4zisAPMSQS61HRwG7CbKhxAM1Z
yUCafpBWg2+UD+MQmmHtUqdO4zEHtCZ26JpiCNcZQy3lDHYgjf2tMVlbdSs5qsNN
3r9DIC+9VaTeJee9Dn606+xr5orBZMnuuBFKgE0aHKeUSgofAS27tJ7jwU8CAu5d
jgjLt5w2eEZgGw/si9K37xwzu6yOiWPGk8E9JofWZzjrPPtO3kGcvacRmjwJpS78
He2ulAwg9u4b8cQCdAhr7qPiG4BXEsWxVb01Mfn/8MqgchnWMYshMNcCZDEqFbJl
0kSp2dGvgveYD0/RE2DEE23eYS2d8O7scSfe/sG/+kY4tSoJ2eiufWdud8lARbdx
lwEiWg8LXgk+MI9Z6aK/Aj/MLRgXMYiNoYuEAlTFfU7mtfnRnv3HqPEZxaS7RCSL
w92OJpnvfywxy8mBlwhFHyCeVrRXprq3fNDAuw9dMT+/e6UDHy19CrtPcCJ9VSb+
QPWbvZpbgFYS7tZbnsD2JZgveBsK8TEECdWPCJ/yF1JxZiXYsSZddk3ZqMTITTnE
gFiYH+7qM6mqkfd8bpqwK+VoX4k6qd3Jg6GjH+PWshg=
`protect END_PROTECTED
