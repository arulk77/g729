`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abJjHS9uMa3VXDs8E2Kh8LLoqHNjgndqZ01XXfWJ1g8S
oSamWtjsy44bOQ34Vo+aJ2OB36gyRCd5KvoSgDBUwhwM3LBZl0CMq0dIf0Nwosez
3Jqk33uFBV6d9WYxuPIE0K1f9di42raZ4ZvryGXUvQjRbDSFbyM14mkvoafjyaA0
2Np/exwIXqiBgiPtBUMyXHJXhvxh24KUnjHeePco0WpqZ7aIvbcO4asIHJyLiskZ
XSv89XrWc30PKgtCdh23KOzbL0CKZJOG9CbZwm78T2AIzZOcCSdjaODjxlyjFY8P
wQTzp5MKkWhHXjeS0yIag7xbWTMfqwxkwBLbEqWs6eMIQBYhuJshxD0kBhemDno0
`protect END_PROTECTED
