`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40NWkWYNi+s5zKwyBehf3bEwGSo/zC0r5/BagzaIADZY
Q91bnRBbBZtJhg2dVdOYgo9D7rHN9xcj0dvqkXI1OR55u4meLrTWEi0NLSskI1KU
v890bswfzwrzFy9e3xXvpvU03dHTDdEPzhnZM5nHOfr7mzRxQqP+yXmHhhvTSKyM
R1RnDqHa06PbP4oG01ctujnpCj69AS1pulncyTIxw/o=
`protect END_PROTECTED
