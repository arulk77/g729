`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zIVAs3SH6ddOnB8VAe2eSs+lG7BAbfPvYOs1VfgNotE
kiLw45KU5rIz2ILMIsFxzFxw2rkuVY9e1sCh3d+87bROds0vCvnwrtrqmDmWwqg7
yBQqyyggJgNRmHpc8XXdgM6sSZuiKxjDNM7eW2KnNY0LqGNlQjj6IiWGXT0H0xdg
1n5id32qcLtNlmntZ2FLcxIljR6Xu0SRxNqQSqUwQgrP+VYunowpkV2CbEw6Y7oh
iB3IlvwJH3UAasSGPIOZyb+I2fkFO8i8UHPLXQkV4bI64dY4WUAd4cqQKWFTlSSR
kFP0L2fBJbhzDbKTY9IhDrfasL4GklmRDUvbWh0NWZWt+IEvzVhNkPYeLeoBBKzh
wDeSv6sdz4xSCahen4iBEQ==
`protect END_PROTECTED
