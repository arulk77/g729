`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44djIfr9r/NJWGNjVbZDA3Ee4dWNjtVOCzC1imkrOMVF
C9BFhSRtaSgX8DTmxvfEvVreBVehMIDgMoDJsRXi3YwnOntsNfNkwvOR5F+rKABe
j7+kFZofJbL4N+Ei92sidy4FOEYocEUXp5YmL9O5XEn14Dn8L+hPPFhzwIV02Oob
F5g6xO51qWmxDUQvG06Lo/fNSplsz0y49iog2JGGitFk8jzj+gvaUD2AIa8jZgyw
XbaF3IFqL5nA1DVPAir5EPNkHMhcmCYfyXjyh1oHQs9f1kUW4faZIghyJEckk+cT
XkAqfLn/7dsNyj9B+kOLIA==
`protect END_PROTECTED
