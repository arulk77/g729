`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAS4zC3+ZJ7K0C4kL65miM9X49/ioQp2zGxQnLdIdbMG
p+rZ7g48qzv3/JVkKf+nLy2+c/u5IncoMDnjMtcrH2RM1KrFazbhvNzUIdMqbt+o
aVdkjr0b6W4R8Q1a9ZWbWX7zBGYpgQ6MzXU840IhwyEOjxW0NvbRkRHTufZzG+od
g4gl0lnm6HwMkr+owHcZsomQCKdOrBosyZJH/VtBcAqygBfv0FjLz/O0jR31uLnH
65cL75XBKd/780rPxjB7igotussy85fkZEIBUD96AWaOcIlvBj1wLIayfSmoo45O
`protect END_PROTECTED
