`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePhMrlMhXU9CRRZ6j3bcsutLqeTpPrbEyDx5RrUQm8+V
GLqLZt6DSQG3+6HkpgO6n0VGaxSpAmA4BTTJS9iwihnbAbkiiB5MNRBESDUsupol
aptyqrs9cPy9PQxCMHeSaZ1WF9D2I0nsR0hep35RfKIrR771peHzZNXD9R+seIwb
VeIxlkGlFdWh6gF1+9r1wHNggi4ExvNEXR/hjspLDhAsZOexnbCDIdPR07y47klv
vUfxl/qjkXNuMP5DOzKMtfmlNKc5dihxsc1CgD9ONg6n5pkoK+Dsrm2FMiu1tvuI
xjmtNMt564HYor5DSAFqx/9M4gvvLgenGam81eJ6C4FplZXATQ1BwNcC9EZwOIra
ZBVMGaWbm6YVuKUUEf/og0vUbUzTjRTS4KjiFaqyCSDayKKrxjHYfbDCqkT6TmBw
`protect END_PROTECTED
