`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKGqeIqWuE9U34WOd+9oHGRa2VRWPqwh/exTQhSut7l+
YwdFgv+XJy6kq1CgN+LHoLnq7nAJ4OYxu0tkyKeIKQLWgWTXSTSbt0E4AlCYj6CM
t94uicLfNfgZam0liUXNj1Ll9Ai3HlNgEfve6oa32ExmfT8YG3/iqNFiDkEz/ZXL
d+dp9OyE334l2TtGZyCxm6xlDaQbdNLMSIsLS0QKsmcKZM//KCrMmTa9grWHf/jh
`protect END_PROTECTED
