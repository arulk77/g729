`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4wj5bNus2kQRQ4JVE6MbHc10bQoolthnqM3MrOxFHETT1VfNsOrQMl6DRCfhO5t2
HrlEmlkZ6cB5I1viVGmIhHXcZxRK0KgThsK8sFdlQacf0hEUcEFEuglg6jLgGhzq
UeMiREfTi/O2DY2LPXe0E/Dso7wj8dAPtK3rx6rSWgr0JNyXZ4VM4VZDXKQX3Qmg
NqdH50m6/qiheEEskBGpgoIBeG0HS8G/raqsZO5NoF77WYY/Cv2Qe/q/MyNJ32o2
Mpwni717hyYkABN7OF5dyUVkLHkei6CTyPiOZxWrCVo=
`protect END_PROTECTED
