`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQspSM4KDPifbiuNX1S39MaIa1gFx48TE3NYk2cNR8SE
OSR7R3ZanmMRiC9eMRUqGijA1qvPYE+uYRYM19OgWDv7KgvbojvsYh5QGuMx2rVT
9C3ITpEDaL/2EkguCbqzgjH1bkn3bw3hJfmhmu2Z+xUXrTq67ldpB9zWn9Nia3qy
xGr65ERkqcrJ/Oq5RbY5e2oHJNytWC8ACJAQXSRiCF1b/+r6xqNsvmGZsNyEbvNT
ZIycuGzfAUrzF7myzcghKNR00ycdl94MDWvhLYUIOOipIU31bMcERuCszHl3rCOT
Yx1e+nDqCjt4GHRY0RgwM55FwzcL24OPUWq0vmam5tw80BG6ixD78KH0yv8de3pa
gAqlnh23hEQz0FeioqAAhl+4xCzRA2r4dK2IDqJJyv+MYmpIobbvVJn5AzkwBjEN
EMH5fAJcVnL5mqx2oTlZvZvS+nDukyzqdycXhuuhUJW+DPw4zq/2hQy995rWaUJq
pZ9WvOTRuD/+P7fpSNQUiNQXylwTh3N8bHbHuRGSY08NwnOJt+/SpYGJOnb/5tud
2H8nqnQ1jSjVIUHDy/B+/9tjFHhHu+Cs/Zp/GjCcmlKfHgoaCSBktmyZEmdA5KPT
fLJ6ljDTcPUSTMfjaGK93pXjIl4BK7Rhh1gKqgVqzL5Fgb1/8wihHz+FEcnjoTU9
mlI5HwVHRWpUSqJS0ixwP6ERJYSaG76/kqqsq20kv+KKsvPaZJ+wzwV2OBULTzjV
B/PoXcnBnEZBH+GKWD+PRM1Ip3FaisrLlv7lYC8tkXR1t0JRwB6DNiJaA1chSg9z
CPJsFHZ4fa98r5PXC6DrmeXyfVdmcN2qOFX8ABRF+tbM76R6ZM0s1fv6wQzzGF3i
Fc1OjJ53SptQ9BuKLBxhOGd0VRBY4m9hrCpaIE2KQL0lEnJJuPZ/MWdYyV2N0lux
xqgRXrHRvdJBobJr29WIJo2rdR4brqKVSHin7hX85gt4rQRBBID1iHN8LUOZ3qFq
x5HNraHlR1NrGTZr5FY2raLV/s3N5D1KP7us2mSfJN0YVuFQ3zzknn42DkZ2HluG
kxj758BcoTm81nTrzwTg+Q1yrj8mff1z+u/FjL29RxGZ5ye5opD41WjrHfdrhVvg
OpWNuj0LLWhbhcfA4OJlAp9+HCAt8053gHsTuLy/ORYhWwV+LqUzTCBATYO9uS7j
8gLs1HHQuxM9ALC4rvXi0c1FpDFC8KWVyJo+oKTsdvHX/BIF8SbgkKtJfpq7Fhrp
ctPbJndC83x2lhz9g0k2vGuw47UAjv1UMYOHs3pyIIz7LbTEMTGGz5gpT3+i7nNJ
Z5MfngSMIflvMPk5CcwfqauaOF+DTzv+eUBJrkMpX3iUh3txPCnG/ppONrhCnUud
45ih55663xPF3vJU7ijK5EjrhVYV27sfiRXVaRdV+LbpI8OiV6yM3BXCk2mBci5d
IXclgTsMPwIipY5F/juFLCQORTy6qZMnlO6me+6vwLkIuS9VK/LMnKGHUhDoAr+g
3/G4DoTYguk3J8BWUTZhnBg1lfWBdUcVy0Rps0R1d+/lXz9SDc/AiH5WiLFln0En
z6VqEMkTD6M6dKKNdPnUhNtjrCDXmDsWJziuWI2qT2qWnqZLj9xIeS/EBU2GlhSI
/HL5nQqpKyDl/OU4w7NY8cl1JEDSmdF1I+4Kqalz3DMSUFf4+cgX3tn5Jkqf+j7D
pwd/JjJZnG4RCSk/+cAotG9utdI9d6ERczNtlABy3ORoPqx/gVcCRPwREUaEU0hx
MaIoWunKMjl+8MUZTN4LXWsKdtlbvgGuiw26i8GyEftY0O/CzCg/z2OnSrLRE2K2
NIG7bukUEv9i0KUnMiW2UjVeJpkCvOi9+5gQHmfVHY+NwhLc2AHQcMBueL0X3/lj
GH9igEJ+7QdZCj5ksi5/RqczxU4e9vuUaweliu4JtyZJC3RoDXmbeNm1nekIIZoi
ahSNzZ/nxxrenjgA7PurcuMMJMMGwGwaIvAI6n+qXSFgj3wiRrRfdkibcWjdKVes
f72mMaOLApzTOzy0isMp8PxKgfGSC23ftmyVpxPUBMjITqCkILFHhwhLw3LhRHHr
WfOA1aF0Cb4uJZW5wCowENcmkh+R014ToJhwb4W2ATWswuZNQlD/3TzEVMxenSR0
nAnPGWhxlddbV897BLMv0LXdagrGFuYeM3HEBUCkMameOHp5auucnQ0LDELckpHy
NsRIbbAgO72L9HcnNLKrBsdhDF85aDV4Xmh2OY8aB4gbu4S1k+fuqTchmoaBM/D8
/aHeN9TRbrX8I0he35W/MthO+69SpaB+V4q/JJoeZbT2y9hhW49bjOA53I62PrTL
AIrTaDG4TxnptIV7GZ9IWhie7SnTrgb4Y0y6jzdoZ2xlsZnfg9/4ENTSX5IBvGzp
zGNXofI1wFifsySVGlaYtj2mxVolROJ6PMjInmuYc85Pf2LLZIh3s6+c7GICdTWv
4UeRiavKEVidgke0MRu5puTKVCOFt2F4910jkz6QC2wFyh4r7VZWlGCc1bRPbMdI
ZFQffx6gs9h4Y9aP9cm2DYpUiJrAla4yx8HG3stU/gTVTf08Tbly1u6OLQwANYGw
7M7YkWax975bs5Mlpmvi3UMWW8uzixPN7LMRvP0eG5ofG+waEsgy0ylsC2JUGYIi
n1G3nAJx7b5PT8A37pkWfybIx7Xeq3EwkYDA33wcrCfsuqbi3KOZ1FLjA21NgRe1
Z+ybjFsOfpql01fOzD8J7BBoPXIJuOMn9lRsl9mri/abP2c4BE8rqkcEZIDpVlPE
RjvD7PvgTDLftjrZTRdngLF4DalU+ct7BYsL2WIeTdrurQZV9jlzFUO2bxVsaWoI
+cmG9VlGh/XlOH09g9Tm/hjDJh8yOsX2YWjYyo/BLk02MQRL6Iard5At8zXyN/+8
qycPk+zu6stKasByZnoOqSy011w0Dz94Gx1iliCYykO7bIKu7hj4bhi+wM2bzuev
0nR/HM64QQNC/82SXOY493IHlcdCAzwniRBc9iRM9UBdV+HtvNUmrmDwiA2jNFZz
wlYV86IdzZOnnVxDH160W2yc5VrRq5eiX9ruMJnpx/nnDctchJuABJbFVbo2DADZ
PKvZkbmxxQcV4HiTgW+4aBPHuDb8rJKBNljuzPv1x0glugXolJqCoqCsLaz2pwEN
VTPTQMIvlacqihxxlS/vDDqIipeYB0EaXLWlq6VP013VpPQtOnSn9jpWeBQidZxL
W3uGVrRKGcq4WH82MBmvenQeta8AVQSOMwy62iF2wX2FYxck2IqZIYhtxGhz2gT0
ySN354e5gsNWIvb56xSVITDb74IsRWKu7AaLetGM+rdtmudbjYft6xCsPlECv6Aa
Ow92qa0S5uN2CFxSd0DZIJSjHe2MnGXOpnPs562PdNYmKK55EK9NsfFGfaSdJEJ9
rOlaxGHCeAeJGbbh0lB1SGkAJRtrATndKESzFSWep22YSmIPN41TOWLfDoVaHuXW
X9STYKyn55GMi2CagjzEmepUds/lX9oQn9QoMoWLdTNzq1cHkYgfpAVbzkJmGzbp
1KP3q/1krOnyBEl5z41C9jDLUbbi5IiOQAQLps5Ij5M9tMFcKu8pBdYHCoJcC0IH
+8rlcZAEG0rbXYHZMJ5IJDkvnIx1B2W49QEP99qzkIrVNTS0e937bb2ODtsL5Dl+
r4Tp2klIrZf7cOrNAkxbn5jVzR+sRS9HR+Wh2h9YZRwOpOqEmrucXrFPhUyzXO3j
ALrjAY2wWDxP0h7v+26NiGDfMdgQ0xXlAhk7/G40WlIj4RqRf/2JGAQpwyfgZ/Iw
87QVk+hVWD67tYmhy8ddCOi8h1xbwl1hpai/KZHqXSa4JVuUG3XGf46j3aMyfCAf
dnZlGcM2H/H5Qxa8Dsy0QBB0FOd+HBKF+UDcE7c7ZkEcmzIuoiHaZHo5E15b4x4v
H3DXv2jvzmYJ8VjF5mEtzGogdMvtLViun/DATULTNcnQVl2JVon3/QQ/8l49bxca
HOBvGCDcsuKpuJKyjFx5fwCoAIyLO0US/Pu/LWmnb7v1lNo7ORedl9yBBNa1FqK4
PymrVfxmRLVPdQRWKHg0sm8xM5a4068Ikt2kpReM8fu/1OW3lu4YyJjEPt5kRoR8
JfI5ZY3qzVZOFC9knVRzsTjxPL1ZUfT1TaIKKd//Xpn90PA5lHZ/VK3lGGSBRt+M
bLB3DPfGnj/cqumglKYmGhIzhnyVelOIhLab0LW5vgXK9HsAJBHmrQP1nfB7aXWN
8YalyaYla7prbvp5xoA9tAerHtUCfBQOHv0Sb25MUOs8axdfr+1N21E/Maxvmt8z
btMMu/IdAznOPKk8OR5fhZ1eP+D7q1mYqnoCioj1hauSRtU/RmVdUcRUnXJCnTmP
tEFnh3uvi8HfQpp8AQbzK60acdcChWRbtZyD4tTzer6NeeniivLlyPScFSeh/Rt4
EcIIUJTpxkQe9rGQylfy/ekMPZQ5CEjq1J/SGO8yzrsbDXzZHoA1VfIcNh0i2Dzw
2Q9r3tIJ2ZPVz6NLz0dGIPXcUciuCy3JKep0y5nz0Xu2/reVU7XO6lJ3oJf1M7t6
lW11PxeME7uRbS31M40+SakBeN8YcGKZ24dmwHSywpA/iWxsbZzS05Zen2cdSywZ
Npi/c+GxsUWd46kPY3UeiMo/kZK44nkgkr0VdwP+8+YTTU1K9psfAdvkWo8AF2/r
COMIcjjwYjMdzDYbTrwDXdeGrwM6FDE5jB4Z0Xvc9InrbYRdT0D2SmU1iR5V1brK
S2DGUQjXwdU1ffKl0b3gbRufeuNjCYSpE0QbE1NgGKfHJ8j1ZgzQO9lhy+5R3UsL
ZZjUteibtYqaAdj8XSS/1eeVJ498sHKN1cEBzw3dHd7MEWGEFqmItzM1A5bBxE+m
SgPqOp6GAGT30o/6sGLdk+PZ/l1SAk1s0PbXOTrCIy2HCOAbEpXLDy0inZvefHpH
Aa1rMXFWghYDnA2WIc6N5RkIXMDCe4aJVwMA8BYm54g0BMCnG3AFFtracsST0g2s
Y3SDdgm5K0Qf/jWhtqBihxkah+NdoHHdBfLtUqYoXz3yJRyN76lOycWj10xY0wPE
kYNjhCXk2PGfx33Ur2VcEe9LHOwLo5J34gNIkk8KdSaZXFiACpdvX2VP+oeV+3ag
ddrCybRzorowZtQmlbsVOsZ+xtCaN8p2fLenQn6VeHqZ7uslQ+gMOgFqG3ZlmJ3/
MhAdGJ6lfHrQQNHuJ6R284TlRRItz5NHGr/0hbc8D9qSRJu3QryFobVeTSFJchQE
P6lbFdgvlschOkImThJRk8YhHy+fNV4SyjUVEmnYbLAV477XrijNyUUHd7ALHhUz
ssZa5IrQtMeF2Kvo/oXIQLU+82tPiM+b12dr89VPhtEhbB4/s8FosiO+9tGjx4Tr
9su/mm99ZCekS2/8Rkej/BhasP5vmjKxSz2gnBRINjlaTc4FF9nPdnfdOG4LeEro
r60JSEgeB4gkmtZFhzqpsw8jcakwyG/RtbvVuh9+Kbz25uQhafLOyq6hnKO7J75i
rrPTEPh6oiru/A43y+fVbrZ21bHMNf/ay21TTA7/OjOfEyqM/v/qJz7Htnr9OIy3
evB2QiUiPljlo8yCZN9MdddIlxRBnPleM2qlSQT8MAPaLKj++kWaqP5pef+l67o0
wTEZmo4Vj2NhOiRBzXNvyERw0wo5dQ73m1IQ8BCqY95WKA7p/LRNiBowfFYh5fk4
r5kv7BqtAApVpT9afbLJWqiQY26VA9cP8sAfxIty9a1+7BMhR62QEx/iKBf+m+X9
GOOo4zmiwTqGgpPHgX227yP+LGl2+FTXgA6S8tA4rkKqWX3ZplwWBik0zP/+QMe3
S082nz3X3vn7o9eDm/ohZpLt7c80i+H6F0QqLuqf0cPa64XVtHLd0KIccxlnT12a
+SZn08DnQHRrTJ/ofPGygP018RwVwvjGHsDae0mZ/iuaqaNmFkVZiyTWiZ3Hgkrp
sJQvLI3FGugpAfDeTA7iaAMQHK7eznshbvQUJpHnzQZsnTzN0udBkMdwiT395OBz
j91/i0A/G6MnIBDRW6A2htWLQ+N+oeC0ZNDadvDAwzqgEI+zqvxFwXcC8zgB4Uwi
AXBAoCqajoiOCPlIKS79Y9U8351BeXZD1qZ4PkgQfo8SIQwgcsu34cuGsmZHWTjg
Q1gClwTJjSRi7TCIofk3jWA19/ZZ+jY9VojpHEF357IfK01WMJus8Fe8XYtMdYu2
CtcHMmQFit3Ltyr9sVkBf50yMsTegR8kNk4PosvKtn5uV57qFpf8RyBX93MNZL/m
BbEAm95/oewXq6YmDua/MPyKz9SSrsNYtZDtQNVRwyU=
`protect END_PROTECTED
