`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C38BeevDBnBGK6Yed0KyZSAl66YQd5Ii+JVxkrQO3dkV
LCsGdWC8cIzmZCmsE0SvA11AJ8uKqVBIA1JClwaE2XGt7SYhahKi0t/ZGRr7JnOs
GpzUGYUFEMHwR5XTFg7PLm0h3QFf7LCJd+ug3hgcbF4sS7CeDqxm+PU0zuCXO/5M
ukdQkkw6sw68TLwanNyWwtllUrGNsUv9Ob9rFseuzn0UM+XcBe3a2sU9UR05tyCl
r1iYcSaJjehzJ0NMH4XKDE2gjozNwvJsMVWXDAGPGvS7tjaBsj5o16ujn1xkaHY5
pbZPQ1JvbhsSZ/wNyh7sVE6zek+ZLztb8bm1b22dmCyhRg6iVFESVPP5V6lceuv9
IJCE6Kc1Pgib/WVbpmyPxuDlauf1n5w3atM5JQKvVxsgnHbFYgiLrsu6PkvWQs/i
Ttt5U3sMms1kAqyUQ+6t9ZP3OW+qM3ugntKR8TQSdBeVp7t8/VX64hrriSiCpKGI
Vbf0kg23K6/wiYWw2/4nqjVcjng5tPFd0ws4vWgrMqkGEs8qidYT6XqfXEn1eRhB
gGAM+rhUAoV20rV/ngH737v/BcZa/17/1/zjLiOEBPY6Nv9iiHHEVqNpuxN1CpFO
Ln+pMytD+k4vC2R5xffV73754izEQngwkgwnurcCt60HbgrQ2pDL8YcY7lWEftvX
eNERp2sYRXmksqvb1Es6Prn9xgcgNz4qeHdvQoGpJH9QfMDny6ZcuJ1siSln/xcb
r03cvRQ8nto0XgcK88evOyVZBIFZchmeI/IR1TXDPR0prBW69UkH6rRl9RF3lZ3Z
nAdUelIZ/3KnK7JFhZ0ulA==
`protect END_PROTECTED
