`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0LASWtQbFi2Ws4YfJkshDWfteXmTQAKpcpTl/KoUskO
EMwtPerFyiCBK/YrUYi9C8SWLdyzNRpCxZpFF9qroIbY+T4HoE/xhXXYGw07izj6
RJtjV399oXIBOoH/uuT9lbxE4uvjKivAX4hZaEeoqnofKsFP7tzzCtzc8+/nQvPh
IcLkGOEC9IVamqo8O47tpzppIf7c5oXLRyG66hdRRxlb9GhewQpr5GIbIKc2EkPB
5DmTslILPZyBsjehpuJnFG3Jovj928JXH4cjMo1Bc5Swd44NzrAlJGhU2boysDe0
1RMBzO50SBAq9GklfcueM+J3dR36XqK3OOerkK5VfbvVIrOPdoICc+iKRjHR9XJl
0pqKx5a9NLznHseo7eQF9HsUwQNTWYiqJa9uKjOHvJTpYOgCT2ryLlFoRf6W/Lqs
km2euAEHT1IsKO4RkBp3BiLz1XSMp8x8RDSJ/+q4U3TnxsL9fqwbC1i9yHtAV537
jRpGQ+rDYeJGKuRrq5IFmCtkpNUp+Ozd+3lj9yOxsELoUwj0HjOOTo2Hok+3hDtF
gkoZF5RErLl8agdvd2e7FsOSpIWvYZomcmFQgz64X5Tx/yF16IyuC2c2qCykVyiQ
r33PR/xhdxxJEek64Gl0791xJLM6WPQPtt76ouWQzgPuHXXq3So7nM3WdouwYnsz
AO/fnFsSPfuErwI0zTqg6PpkeoqYv8cX285Grk8KYKvovWHPY6OPEgsTrcCLyODE
huIV6tfH66IP5b1U8JRex/R5GjM0wTR1p4jGjvwu/NRafuMJ3x5aYrHBcXrjCT/u
C4HrmkcJ4Xn1p1zoz84vTb0QZnh+bbUc/94mZTHf7JEGH3vxL1ceUFwOVNmSFYF4
coifYSw9xoy30XIYOyE455wOfVfH2RTM5XawqWTmR/V+U+MCIGgXluPr6EVSrxzC
XEzgrtE5SIyVxbdIYxyIDEKLJN2EUwiaaK/Pkc+szw/e1Bw+1yLVb3KYva5hNQhX
ixnfrgfvQIJbMCCRq+jl/tacurpk16e0r9PLd8Xwb1YGtkIk1UKwGkdPBu/NanOt
qhvN5+weCIgrwsIGgC0hxKfV92MfgCy+srfwKuLrSgukYWsp4GVO4enOn3PmmfqY
Xlmdx3qAKwdpMk+lK637fg==
`protect END_PROTECTED
