`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49gWe2DdsAuFWqGc0yIxdNMn6iZHvvkZ8DcsWwwIrE1Q
lSgBj84wSc6rY5eY9ke6VYdm2f3LAUniv7TP8acUmifPOfb8ZZ0zR2pDYe+zBAIr
H4XgLCj76T9CZePKO72KdAILBMItGULFUMLRtdU73zlFfNGfK9G/7gzSaE5I/M/s
CsjFetyqLtHIQLtf/+9ZZLuacXq2FykuuwGUs+eIo2/K85qqAwhS3xwAFmVh8kYc
TOQufSNsQ+mbnI94GhJuk8X8RpA2AMhMYGRU2jFlxXqF9ruDaX0Y3c8XjRN9Bd49
xl2M6zBDeJ5KwW4tuw5s+g==
`protect END_PROTECTED
