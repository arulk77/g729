`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMNuFtOCjbxeF0DZ1JxScMAmdjB0WXEof81I+N4Yxj+O
DCx/OtTvO05ZDyvsrm2tUaxAYJKr7Z3SOdK9ttwBTQC/9wQ+PC0MDwxDJDExwzOE
n12CHwayKeHOf58RIYsIAAZbbg7meDr7j220MxE7aoaoxIfBmDL22krZ6K18VY9u
ER7QZIzN61PrEwDsI0PWxQ+VjHsM8L3iMQZy/p9cBNMuYaAIaVkmHaUeJlQK8geP
AUS+wxfvmo5o7m5p7WjieCH6wIMnQDBU9lZhg2EoS2g=
`protect END_PROTECTED
