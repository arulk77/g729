`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BMZlZ3qDES+bc//XUePh72cK6OK2RQyH6Yem4MvHrBKDqLKZhhVwuuT+oohjZNWx
g951KuLQNXTozBKyggcYZ3eUPCAz/+Ihx6eDqJWURpoMl8/wrAoKxh9Ao5Yt94Ml
oUSYJeiu7Qna0D0FwMQKjJ/Tvu/3dWd0LW3E4eLddfPVK5CKpbE3SoqAepBm2qc6
5aLn71YNoDjRFga6uARVF2u33PkL0YFXemNtKh4yAgvq4yhx0sXVYyf/ez4Bt5OX
zSflGjV0BnjT3fkYUf7XBMrP9rDKYF7pCNStigrhUis=
`protect END_PROTECTED
