`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKxlW2R0ddw81ibTF5fpb9o0zzPCNoT4NqP3aKoyCeNy
9EC09srNbb1V5q5/5aDinFrnriKeOBrw5oA415pMzbv6WOI8S4qCtFdYWfKN8b/h
uYivA8JM4gx1MEjIwBMsbPWFFtz/Tx0tHQWJQy4S4Gxv7LUkTtxP7jOjNDshdt6O
vzf/Be6isa6tyVX8Je7hJH2deIGouPOTHNc0jxdVXkdHkDUGi8lHaaI98So5xGEe
y/SmKgcmmf8yWkh9av2g5NSVAxEiopHoqJktD2qqsHrU0aK32Pe5KwNQyPmOq/FV
pftI68AnAmr971RJTidphgFrrUIoU2NskQtWZrulbKeQGjPRk6kf8P5AvEVFbZ7P
XbhQvnB4yjVado4YpPQoJv7fintDCNueSAcxqGDU0FeI55Z7khnuor317CBVg7iE
/92xJNQzl5yTDyshN2wzudQ0d34jBB5/GdH0r4zSoAiuqFxHp3Zj7z+/meK+1i5V
`protect END_PROTECTED
