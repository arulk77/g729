`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLkjfAHdrNhQnFpS66IhTyVs+D9CZ6KOxPrDJKI7LXUWg4
qVG7Bk6fjmKDGZHSr9WHN3DUXxF2FATMtDyU3g4eML961nfjKDAsc3agU5zKTEYo
1fVcO7nwBcIXLKYD6HT4TqYoRxXQdKVRnMdO0w/8to1ohDcn/mWGrFCSeG67IS54
5KSJaUlxBp3WE3p7m4FZTBcXrJ/8k1keXRtNsbWep3e42ykjpTuKiUUNVKjNfr9x
yrFR2JHV322KA1zRMwgleRMIZyWVqofsyHh/Xg01D8Adhddh7mb+PJ5OHpsLLj0L
`protect END_PROTECTED
