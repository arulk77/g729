`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOshMJoolgNG+47xHytzvBNd++IiSgDn6c9m0oc6YvLh
WeIDm2kdvAI4Iki1C59FEmu7BuSGaTE7SddiBH4bFoT9eyPa7xFE95tK0EUWql9e
AvuBViUjCwc6BAvJ9oOLlOvBMpwpIACfrVrS8jhM200qz6UxI7P1dZsPI62pcOav
mvFVAOr9gLW8Osa1N/Sqc2aub0FImlVL+WVzYYDBkq+Q9pwTKH24loPg8c9aUGqJ
gdyfEuvJhnKqp4SZJQUYES2xqSiIujke8Rf1MN3Bt8ffHYQR7x/m+5j4QKEV3ovB
g10xAQgAN02NkL8i/nKeBVLBw6e1CcT4U+mCQ4r2Aac7j+cjiE/dSwjRXHZqXXlp
kd/qc8wTraSDlxWaIivXWxhVRG1EKPt08V6HuH6WVB0R36XxoMUV2s4Bs62mF6uN
baVscpFMtexB9aebDf0InA/+GLbflPhiU0tnoAA84swafYw0WaDyVuUUp6l/XTDz
`protect END_PROTECTED
