`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIhAHUuBOgwSbQ7b49Udo9MF19l/dBaRd4/EH6qTzNfj
R4H0vvUKHQ0tr99OYmrb87+NJshEfXPc4d/5rlCWWEudsFzPZvUQ4xTuH1i1e+Lv
DMp5llI2O2iISO89edmY9esksi/urj/63nSrO3dZ7xjwbiLkZg+XhGzHCxRMpFwM
UCvVri97mcT1t22Rxmsn6EPzZ0G7mrlkQ5CxkwOwUcg0B+LOkIvnSNdWmudmck6Z
YpdjnHWGriBotaC6L/ecey57D0nO3NzQK0m8w5YQaUOtVhW26DfRDGrmfIRR3eZ1
42R9lPcGqIZKg7dpK8L4bq6I6TMNMCjD5iJCC7mNfGNCD1kaxWf3Lje/jzS3otay
LUCEv7x4u+AKWBVSuTpENPzSJhgJ7z79oPyXMn5t66BbuOLdKXg6Tuh/7HzRKBcg
gmoYyxuEvNA0t7/+MwpF6oCVvORMpSyK4mgFZOy/cxHn3n0i1T4y0b9XwnMYws+z
oSCc1tMpYV+/xVvt8sFk4TL4d5nz76SP43TyxVz0k8p34maSBgN2uXZY1h+be1pr
5iaof+2oMWv386Cdpn8U7Kb0gz1tLI3LvoXqDA8VNo5/7PPuLSQ7fDDDQMfr0LVt
bXsownTDQ9hVkBvy6GlWf6IcPGgPbhdJF6fr625kp7jZ4LCJ3syQE9zxlfte74WU
`protect END_PROTECTED
