`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GjaMtuhxff4B13ZrMWBjmd5n9bAz2Df09I4FyjDwVjEkimN1X9lsxh4icECNhuvm
Bly/rDA1c+R/3n7G91cX2vJHNEQR7O9UE5wbyJvDucPgQN4RSFHg55NV757h8YNg
A4oUIPcPPM3n1qnV+fBnCn7C5eGd2ysf8vOLI/tVX7sQ8s96tprR5Lrhw/bGBZWU
9X2e7lGFN1R1cS5gCaa0qeG2+JQgFhFBh6rKqgiOGCM0KYIWQMdEy0OL9QGr9ZY8
yVnvwi2Ot35Uwo7N7tdg5PcFd48QwvNf83iIDHx6/7GJ5psmdnNR5Gpp9NPruhC3
kBrtfN1rmn+sLczECv1EVgt/mUVFW4kDghi0HNG1HzDJ9MOaZBB81JUrXGN7H/iJ
4wgKrMT0NRC+Wl3JOoH9MKLyvQ2DmQI1mQXKDf6gfQ+W4sBfJmeRn8dRHLjEGISa
o0Y5dijcYc9AHkFXhvDvRxRb2a1K/87CGQqSKWEdn7C1rw2kFwaWROax2VoQAwXP
CtieMWy5oCzG8+pB+TDaDRDGJLSy36ytNMP6w9uGnJrvz7tNMG8bb/yaZQfxTbzM
zQ76+oTPsSkf4k0SU5r0v3kg/AniZXswcGfI1lrn2rsPfPkds/+wZ1bZDmr9DdgB
4cD8tyHvEj6qXRyR891atcH74tSnnXc0CJfh+PF+xjby3MhK6ieUUZiWbWEbORIC
fdwHttbKym1QZi7EtSUA7XouJFucS27GoymsD3dKvX3LXhZ56ZtuLPS/rBuFfUqg
S8o+e3PjMcDoLBFImzwVKwj8XM6aAqPehWOrOCLcdtmr36S3VVT7vZmAeXfpSsTC
i6QJZwW1Uk1Q+/t3yb1aKbJRzwYlNDzylRfgeUT8Ii6XXxRKGQrfiCEtluyUKm5C
OIsqIOmvO/xRUethwErxPDj1Z92siRZx5UvwBQV3kodzNSjtPKNc4D+/WwozNX/B
n9Yw85LCpM7CQSLFc4RfEsAPj9QG/bOzZdYXW7qp7rulH4Pn5s2ghKvUR3lEK4h5
e2DI8eOPZooGD5IwdgStYOKHFUat/MvFuHjVRaD/gfEFBjoR08J7MYE6ko0P3MQH
28vZOh/cxVqDYhEbilusO6znLAnqW1cEkgPB/qzrxPvZ38EvJkp4vAa1KIk0348E
z2IXrdXJgYxoI/J/GuzGxAV2n2Kkp7Wjx2QpV0PIDhivD7FKljdO05MLF42nB9bp
ALf8Bt55VxuPd5/7rKuHLckp7KIPfg2IxQIqKwLuqnucalZfqb8PUJ5hVt7fE3sv
mNE6Azj4Lqlxkhol9P9Z5jisB4hmS9YOp7KBiv2J49GRTOJ5m22D0+cc9hi+V/TJ
ZdYtgB6t0ooO7F3CQbtyp7t7ABxaCuk4XwAvKChAJuo1rxsJJsUJXXKxTxbDVDSX
gjsyraqEP71s+AmVUVQrMcE7eQy/OJbBbbtI/mGAPMQmCj1aTuk0zv8nH7+/yC66
lqr0JJilRbbzDEqLgeADBTFN6dS4c1bON3luSENDoGpzCegleE5ieNZCPIfk926u
oKOCwBqBjNkZmS1JvXJOccaqPdqSCepe+HZNHase9OqhL3grukGXzGA1Jd4eXuDt
oVTloC+KIPxLH+P2ZlvfGxfxe3/WVfkoxrnlcO6GMDvCDmOQl7P21EImc6PdOdG5
n25YRGh18S4dk09GDCWtuFa2tbQ3Hr5d0qVjeSjt0ZKIeTA3gC+gzdz5KHY0E99b
jC9gzW+gH4ts4Gqy2ef3ou83S3Audf/kI+vpRpPaBLkb8NCu6FYxoxeRt92LiqKC
z3xjWDvkQ99UgeWAuB382fMw6UZGNBte4LHN7aJ6eBcq2TEiOiWlS6maBFlrdk49
fSCGmsvF7WNP36PaMbrR9Bz5Z3kMyKJiQaigKa+QAniO0tDzaAw5FpP22QdnYPJD
DTuZ87YUheuL3BOa9SivnShL9l1rG1Zq+Th5grzv3Gfpf2W0j3v1EBpozplkGLHS
Qj/8L/MelUy0SD5pEPGolOlrS+caKHU/juJVG/0hhtNA5CsNdFOMQrbcbrePVTRc
WWXDp7NpWK5ODCc8Nx0A2oQrMs1KN5P6q5L5dULi2q8EBTcVfPoDNOsAI6P1KCBf
+bUskqN9djV5Q8OrHrZsOcdTQBvm7eih3AwvsgQ+KmKqvCMX3iZ862iq8G3Mtm0E
GHLNXVuLXDu7BWPWpX4n50VFR606Ce61D2zzGS/AyW6FrmpYtlGgsV1rac42QOS7
zzfrcevQOio/+H3xUYAFShAEbKDCP4xPyAfPOvUuwvAcUSGsE8QZzPl0S+Y5oDyj
aUcgDuIDZjqmvYx9j4ClJkQKOwdkH3bTMzyvYcPOk+Jplz7EFN1V4ZlWFU35dDLf
cCklaewbLc7JgmdQOJqBNtRoKRm31r9naX/bo5nKREgaFcpJtoR7kz6+M4qlSGdA
wtHNqiRZZcfmj6b6gD/pAG36raAHWB2xsCb0vPU/rQ8VyEH8uWGxA5xBoqH06FAs
V64S+DYioGKhenYFwbyxM+ttziqNc22DgXoi3jhSHpAFybMzoXeHDDseP4lWyjGN
3WKv1YSdiuYDmQiG7IWpRCq/6N9EVs6+9sE9OZPloJ58Be4pmIJ2ypFhyvVQvpmc
wFgai2BmXZT9lEFF15bNbcsbWGmi82Tdwo+zsrZ/BpE3AQp1Ar8sEvDGzETJAea9
3lqazriE0gWkxVAbOESOnc+XnQNav4tRZxMk+JNWHqoMio+Mo9cGx3rn75kJpN5E
wGfOPn9Nf8ynw3pb1l9r546Dsn7Y7YbEFo2SpOW/bl3xd30WIo2Ku+lUK/su29dI
hQuzk4de5FARGXPvIENVXCimk06t6QAy0IHsX4hXZn9WEN3PRX+uWZmSULeZxjjS
imYTW7CIL87cPPJB6Loa+ZZrDNkBizAyRQ1A1d3bgjLxIG2sUFANcudu1lzqiy3H
qgVcvYBJqZ6YLM8fn5+lgG6jb6NnRGN6tdjqFHXpgGzzQGZTfsRcJrtJuTzmMEv1
2rJt96E+0F2QRzzIMh3++/+mCOBEDBVA6yv7fg3elCt1IbXxRkrITWTI8zoDMsbD
yeluZjfziApvjoh5gh8+FrHS7QvMWUiBUlRHw7EU7ilHqVGbx2UfO6/D6JhfnMsR
fNh8ryk9fPlhOqhT9XQ/w42LzVQWpMwNrwInmH1k/T+pmji8yQhWbwy0kY38fHsy
LQ/E6708dXJ3/ax961LyJr0pn1LTD0dYHidbpZlRQ6wLbLUr4PBX1BSp5XZGqWbF
Q4Ps1ypjDUNwqDh32VW3apZkNXsTM3BxnrpTiQGVyIU7OxjpRyM1i8tyNxzGcK5Q
Bc2YvOg3ew/neKKPB6ZlfyRNtT1+Nd2zkk7sQZTzfXAi9hMIRhe+4oqV0NnL2ycX
vsSvYBVQwcgKwTweKNhVhb6Al9L/HPzA1t5aVcqsfIHmNGLuqqRFQ5T0GmEcb88w
xgIoMrjj0vjS9Q8YAytJ528GFZfmfORkzxB80gjbVsj1DU6MGjri+RIWi+0aB199
brOeY9B4wVM8ms3gfsLjCJ4I73K/cNqD8Jlc56COiV/94I+st8bsFuLTrJOyDoQV
Kd6w74gCPmbpeijtoklzTCJRP4zsEbQjRt/ygyXgrIpqHLK5Xz5sBPgQS44WyX4+
JydRDY2CWNy1s4VolJDIxsfwokcP5YpwirfvK+w0U/DmesEF9mFXy3hBTrl82DEn
fYxdbYz+LBdSDIonaF86VHvZOV8cYHOjLHo0vEZODHOB6W4slBfY0xEX03JIqVlZ
ZYgYsFnHCwm4DqgBUsA/Snjr+ROW3QD4j/wyJsUdK4zhOJzo1G8nq3FxHAFQb/yt
LK7OZK2CCf7qNVNnzPYrgZ5I/8efZPLz0aseYnqqR9pErp32UK2iTRScZz6KJ9ic
GvMWv0C/i8gnOuLo+f7uDo3vrL5vkcHVwAuPN+OaZzdMg1+4QaCyQm0KSzTHFAWM
Bi6uQcGyJQ+JzAnCCM6o66SrExc9z641erZBqdsf1LM=
`protect END_PROTECTED
