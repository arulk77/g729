`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TqZxooc+4JcwDd+yL207U2uOJQHoDrxsz4ucWAYTRVpfsM7mMdgMRHX0FYBXR77M
k3g8jh49WL1/YxHp0ib0dEqHSfbqSi5z75SurNIh0wExuDEb8zCu51czUcHFkBgx
hk6HyTKzqaP5bWyQ0L6/EjNxF6IxkJVbUhhItAvK0qcjNlwLP661uh0ITv6ZFuKP
f+pbjDnmPiINDAxhfUCPwP9LBeNsTJto6xrQsFI48cBLy1ZFfDjGeO2Qy0WBaBaL
KrfDJyzoSuUSyCieSHqTl1s4R3g9JB1DRWIaHiksrIK1dmd3tYOkvjYlUuCb2Mo0
mdD5GwKaIw6drgKN02W1igut7rlNAGC4vxKzd1AYRSo=
`protect END_PROTECTED
