`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN6atgwbYutx9+acCbKQjr6tV3lrwVyd+Pc8Ug5FvHsB8
832bOWesdH5UwF2i2YRTD9+sm4oKdsZ9QoAXmQ0yZt7odZqIIdCXRuDVNQjpll7I
lZHQgkZR1aE4FQ7DA/ilz3fXlBtdvNaMUqagS6JByemM5jkqaTTiZrN53q/YtLkY
SyXgxwHMat2IMNQq+WFNmo3nOzkAhobFRIRmePwPS1F/d49fZaopPhg8V17/O4VB
iBYdiqi64wppzqrRjs88KGFTpK+FShSvq/EcDTGc73PchbcHw9IhNmfzK7QDYKvx
u3sk1N+Ec/sAQNhG73ekYSDteNSr/9OPdPWSvDGUbOHNCrPR/grh/LtiRw/f3GmB
NHpDFPtRiqZTKiE5i/L2KhC9s7PnC7e2Ysjns3nTKvvKc8+K6G3hEhno4l8eZnbs
dUj8dixuy3Yh2z/pAPUn4LGKCuDFxRKr9y5OTMDaNkh9nvItBEDKqecZqsH2kG/F
viTxRT/naoA2N1glRcStPBVONmntgWI+i40Q+U/cYP9W2UZg37GZms2lOnLDElh+
BugsYaS4YMynRfAkaYQV8rCgA8PA3/nkVLGtE4qAOURmRc12XQ1dnV5IqlwLsHiD
qqebvgC2HAJIGQ8e07gdL62cYRSyC6ZafIaf8gEzYdjqmw2W+995M65h47JuOU2j
KkBKbP54GwNIuxcAbwi2nlYO7uq6x+Fl6V1s0SQYBuPSAAHdejYadQJF5FdWVAGB
2UteU/FoGlMxRNwoWSMUH47cilnXw/XBDmzVlY1BlN6YF4xyOI3obOLst+m8cCsy
jlK77R/nXlkArJFRv2Hnhe+ioDrr3+RP9H9gH50PhG1Q7ZYZEfJ3XFM1MjBHk38o
4KZF4uq/8bDIKwn6cCYMfsDq34GzpkvVaHIq8LARwrtqQnU3h8IL2AS8QuE+gjIS
2YH3WQNWY96AFaGL7hjrvkZ4DaWpuaq3xj6J48QH1YR10sBBb5bkX+OqVgGKCgoy
V9XaqTs3A4l7DZZlxNP/VvaGVaRkue2Kdors9tYvHDZxI4OnqhybUab+7i/7GrOu
pZ7wSWlq5mPWRh2cCtPopCQiWZ0YB+QHRQ8fpi9lm+N6T7+b0T9X/yom4BnqTxcO
vpAgNE9RFOSSMZQJ4aQtGrCsy+B2/Ets+ND5pR1Kg07rhw5vbNEd+FXIw7tUv2mo
a8RaWkz/qh6VGA22EXWOGIJOywrB6YytqhtqMjh9HfVjLe96Z6xdvv+Jzv3K0aNy
UiLOZSafvWqfhOwJe3Mhe1i0LeJGj/pfmOlZqqTSSxzC5wNhUSK0UYdW6GUUXh+j
a+hKG5Ljy0wIxweYY3wxJByQVcEj7IRC4/xTEygNxiRzPKBtML8nyWlOPQgRQVdO
HfOUzRkSt+brDxmEd9u9g2wSBGTzyVIA6DkuT5qweGJ4MKSKYboqfbSTRalfIFy7
DIVWgWjbBI1RMIpX9TkUUTyZzYruDN++K/vDMm+F+9w2haftLxmFDA/WQf2RQ8OG
p5OFi4vOi/7r1jdVlqwbst1aQc2zUJRHIUEEu8HOinBCUZrWXPO/VUkeqyUQGZDt
U/gWoA0+h30Cl/5iOML53Gvp9YvkV6z1Cj038Kl6xQFScZNTMIf/s7YeZNq9+cfD
ehxdanKwm3irfwcpX35M5s/IbjHgWKR698DkdKBwdXtJEajvna6scopfed1lZPom
T4Q1RNz1ZHjVVZIJrIHgeY1le+ZX3hEq/N4RUAWyHIfEOXfyzm6/oq+wNNUNSh1D
9Dg1vvbchtH95tHOs00acOZ1mdIMPc2VE+qQxunZIiiCoKZcjthrQNx65p/rVmQC
+mg2m/X5i6JfohVrZpM1gq5N96xhLZ/iwwcoflam1HQFgFoiTutuLdSGt+izzoJu
HQhZ1wOidDVJLPGP9m1PRbugVhNjI4R3LYRJHxnh7T1uN2Z6RiQfHTYgDmXRQ7IV
0fZ36BOiYKEwYBK1SG1WrL4xL0/ZpAeVNJFOJ7+u3dxS0cAhyJD3HpUvtTcwIQB2
I8fYw0txRF5UMvLhyPgUO+DwZnsyeCIV2dGcnviclHkUF4/7WNcJmSGrd1hT/nC5
5xWXiJIqiEbFKgxKxiLfI8SnL3lTB/rtizBkz40LbIwjE812l86a71FY204l3mvM
vYv/pXDoKv3oBZvsgYUSZZwSpkmjw2FACjzQix+cI10=
`protect END_PROTECTED
