`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
059b89Z7T5H8nnC1DCS01JCjvxPnkDgQh84KMp6v7nTlAlGrNhnIihTlmURoRmA2
NyIyNLb2c1DMc1kgehsnaHPzBZXBe5NbzCh41Y3rcG9w4kd76I9nzz9Pg8eElToz
`protect END_PROTECTED
