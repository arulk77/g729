`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOtgg7eID0/rm+HL/qGlf7xeVYc0eIeHYXKVi6+BbT3y
trdk2AgfxN04HODvGxMNJ8puSjoBJZb+VvHzke4XEteUcv9gm03Hi52QCsUdURhf
29h3XLg8a4HQOMZIw/GK6sWaOYk8p/c5DAhD8j0GO23SLVkAFn/X8hSpiHGAstI/
7yaGvpzjwy4s7ssANjMqeYahRia6gOcqx8wWqyIi+dRO2ehxW/nWuHUDaIUFNOUw
OiUgTpNs5z1ArmJ6Esw/ianDcTK6Wcp7kxcIOWcMLg70y7RRQarXTD8imhZBBPmJ
Wu7wtBonV8rEqwccnanyPA==
`protect END_PROTECTED
