`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD3Rlc+re87vnshoa/VX0/BuW7WVThT4unUgySxb2xnE
Ac1XFEyj3lemfAxUtdLnjF+arSl6HlHzNEztNhJ2q6Y0CM13AAfNDJIaUJF5qfx2
N6H/GOKpkJhVeHCF+jZuShUkHS/pioimtIqGY5nPbxsjTWmtC2FZkQ9E67Ln6CuL
17CODaGFh5evlSF2NKx3KakZy3aHZo3odDpFj72HNbSBu5R+t8mxD+88Yrn+To7A
2PO7w98c+hHIhyLNWbN+0OzhtyU7UOUEMWsbrzqvf36hO6YJmoEBSbRqK4V0EJj6
2XN6hiMxwfapzALvFh6nPA==
`protect END_PROTECTED
