`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOLz1afBcPYGwDZN2TQe7VvG8fTLQKiLmQx9tOpvLCxJ
qwN6EJ77oJmc+Ntk/4y06uk/6sqF/PIKc+LJW2SJ2K/8WbW5E1MfAz9i1/+OAsif
tFSNRHcILGackluRCssOwLnLl5e+XUnL5YHDZPOjvSsYlYNNec3G9/qLgTA3h6XR
`protect END_PROTECTED
