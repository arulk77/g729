`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG455Tka6nlcfQSwyBDajOPefw5MNKvPah5QhyWkz+BP
74+YO4/5RucTWrV25y98GNSbaLCPlQ64yOoQret7G60HXCQiILvJP2X2EHPfznl1
QDuG4QMzOUmQoAtjFICYaGfPeTBE8J4ovY6n75E+QhSSvZbf28IT0KpazdytU9lj
USnz7VUC8N4C+xyAKL9aRbfd8FY+/6a15awJyVPA3gU=
`protect END_PROTECTED
