`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Bp+19bBP5+hB6U1QSW3XH1ARHqcIqfDd4XopNA9JfPvYV3XAFspWzx2H6cf6WrhJ
OnqhdAs2OrSOTKblW3g/M/Ptou26WcNJ2bQF3EdMQfbQyo1Xh9LK2h7oysudVIpN
wlnRtfM+6+ksB0hxbcXbcxXfCWexqJRqvVelQLQjfhIq9/oopROs5/6p9fw2ZVPJ
HDGRH93fI02amn0MXrGvL6ruDXLAa5BCI0eKi0AIDY3Au34FV6hQZis/zGHN4q8I
1gYJS68bmebgs/zbc9ccobDQ/R7/tsZ8BYH/LLS+qGE=
`protect END_PROTECTED
