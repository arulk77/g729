`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2H0yaIB8j7073ZhO5vjQavYIrfx4/1QDO6ITOLYt/bYQqfReY5RMEFwhLRGXuiiC
+A8DypDyUoKQMT1BHCV2tI9dutw+Ilppqb2E9ftWJ7bGjI9azsAFTZX9s24X/r8U
YmUj3T7N33UtURqPdshDuzZvnAXMSUmTTRIoy0OdbhvfnYhGsCdJWuZ/CSYF4ndu
mDMmZr8QipjM9cY5r4nnywIJcrBpjxYxnI4vidj4PnTjPBvKr3Wotp22o3WCr1RO
+w/Vt8xwvF1LQMoWbHBITx8iaCTqoN40yQCjzedTKuTB5547KiBkh4kjokRZm2VM
p2ZcYH2T/tbczfxRyADeRq9BsQ5qmceadZn/bP8HvP/R2nlR9zlPCD53OyEsaj88
Sj2T+N2BICI24o7dGA8Etr+iwfoun9gOGc9Bq9gbystwOjQFWatT8LgvKmh8s4wg
LxxREaqYY3wG3LkkZTTqCQOsJkV9xqPrCe3J362D7sWyq7avvQ3b16RPerRvLPZk
235Cqk67Ze1BbK/m5WaUFiM2G7GCyMnq1Zhb6jlgyhTubuTOy83+n7Z9RF7Gdt3T
gsazzfds+ChKSNPlHuHVBiQUgL//KIXPx9A6LTnyp9uFdD4XcZ7fbbXLTeVoOLzH
4gxo+HX+mPFlwYyjMqXESQwNi+RfDZSK1CZ3Tz6RwHy/RwoT0BAUmw9/w4PK8w3B
LptZsSUASEnC+/hZBZg6Metu+n1PityWqUCTWaVUCGAsQpJWfEdll5hjMZx1dTmc
Rls8KQMcORpksyqV6k/3kQ==
`protect END_PROTECTED
