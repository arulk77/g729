`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNPSvNgA6WX9byDEnzUOb55wrJmZzR+Pkx8oB4omIbDt
QbGQzjLkuAFvOwXQYfmh0AklKBb8klBAMTwfW6VuNQPlMA0A9+mWj+IQlVtZv3Cl
TLx9ecCDa9zzlcskvPhSIt4Ll5DUc30jeBrZkrEl3ctX22p+nw9/P+76yzkRQTMk
LtqsapGyLit6slhQDmH65PhtUTfAA15EOxu3TUIDjva1bfcqYipmEx0SI4dTS0U8
0HJA0A6RTLslLN0Kr6wS1QlZui57tBMNJbhg5EE6mJzJMJphN06gbBupOKCUSgbP
FR+bJhuap+4vF414AJcrt0F5SBXUUWHwmjweuYEGhVgZ65vBv+60LpyDMtjZmEbT
IZWZyBoMv5R+WXBoDctrNKwxbODaOUIYwq09wVAC3LpkXFAN5Okv8fo3NKEkjNqg
yegcgymM+DoK5eJyMB54QS3CUMdyHopjv9pRsfZHtUFmejvIL85DyMqN1bkpqZt+
QyhxUlrXC1tAUN5ySIy56Tu8+6C1YyZYtiVjYRXBxnSQqcl4IKsu2FOZTEo3Ng3P
UzOHAIpfolu6uRDLxCnA0orU7v4RbiEaq7iwvBxC8WczJGLJdExCxJ/0q4ldpf0G
YBHOZzZri9zG9Z0qrQ/mhJEMHIp4Dwd/exhkWQgW3W9MhjDz1rbNKVIJI4zcB9AH
yfoXyLsSHJormzegdqzaBILNvvq6yRhZxEt/5DfhkQuwIbDbyf6lqw5YE56YT7JU
3IUsxl17eP2S6V4Zl7Snr8lFIlG1w4f8HiJ4kexn9TkfLr8KoSyI+hKFaaMMRH65
YX3Ah6jUm+MxPebTlVA03yrrh7nd5hBjrMvicVD0jOo=
`protect END_PROTECTED
