`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aTWBTgRPW24uqTEmQlgIzcce/RCb9CJeitWuZX+7tN2L
hBwvPEwiIkMEfuh08/dOgGhi9FvE9qG+mYiqTqLvTPoiq+XvatHpyE9XthDO5oax
h0Ln/X/bGxi29wWu6Y6sw9p3IIGptGURd85wuthZ3B+wdbOkdP01TgBFW417y0uc
c96AvBCo5O5/UjV8DxAIhErggj51Bw2GGqL5T9PWqp0b1DaFUb9qlWATDJWhZ4dU
VU1+qGjzIwOoWkwt/+oLwR/ck6cefgw2fvJewim74/0obgAWooLZYmfIGTVfdVN2
/xp3f3yxN+pqeEcMMLVsImiljFJnkRh5fE5RqrhE7uToUKbpHRb2lVN1s2g7ts9y
ZrPiA1Q30Yx7ko1SUvR0ktDQu5C0rzc52mZOIK/I0gMkbluDMgUzM8m3ox84C7r4
vKk0xWxF1Cx+KwoUDLKGM/IB8utDSvjqe9QwL7sx5Z+2NDrvYhbJiXjodLQLu5Zv
ildnVD5nTQrPGEPN+wjgG8uh5fzLtSc6fCX0MJ1PLm23hvCSAS3ctKAoWqbGSAat
Ooq/KieuB9lEbSSVr/Jk1umk7+ZUGNEfjp8J0iXIxrXDioz+V0afCDlF9eS5Tfh7
HJKobsJfMVPVg6ZSwewNzk2RJELzn87XwryWN0edrs0Hiy14C3qqcOzeouR8L0DG
4DW1YHhreo14EPksOJ6rvs8jkYSoY3XtHrwQdc748SoxVsNC+z4ZK9WKE5a+Gyf7
exYW0x4wb5Iz0cCG29XgwM/fvGPvv69MQUIq6R0OE50RCGPhLTI3gH18IyWgmRIY
RM4EjSdI95KTFyLk7OUEXv/NmrPblyU2gnlKnTNEBobgvuB2MS5vgXUPrqzolcr4
Z4j9UirdK5hfCULu0rV3A4DS1cBU/4yTbJakZxoQBimnUSFq71T7zUbW8UAjaSyr
LNOcx0fPWcotgY/8gvjwqxCiXGLXSGoCoY06fH4C/186J3tURh/H7JQlS0OOZInT
Ghj8M1cAUH9OTJJAQ+n+PE+xw66S4XR+/tHHnAp7dsk8l0kfj7wfEawGoxvyX4vJ
Qwx1LQucCqQELxHr07qPF7rPEWn9ur5yPVq/kwE/VoR1t2MEHdeXiFDDTfnF0Szz
tPI4jEw4/GTLiWPHsINGD1J8XZEIQD2cRjZ7kuuSHqAWtXikIKR4w0BJ5mUsDwET
M68sp4se67ulQcgy4ldV1XblvW8d2CzChVCsaUz4rRtT3uG+xaYWDbdGotkubCkr
ta6snIA4Tlxp4V4yRYSGOZlp4a2MPJtQiG1K7aOB+aKABWNJGc/ZFDzOJ+YDgZ9w
W1AnmxcPWAGXR0yW1+HtMKKZfmcT7gnWBVe5SIEMuQH0vhAwb6YIyvkmzQH9rV9k
TJKuy5NM+wqdpmHKlZx3M1AQngh/RQvVDOJnR9/kR4QRSsOWnR0+DCiLyeUH8h5F
b3l28S2r7BSOUK9oSTOTSD7wC8dGjWOJnrGE7nglg/g=
`protect END_PROTECTED
