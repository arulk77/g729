`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42/pfu5Y319oeJY7aeKobhtff5EhwihmwGvJg0ctNHiB
blPtJzIcJQZPy3jMV1j3ffdfL1Mna3KeEEKYJYGf+ZgoqEkB81DAEY99YOHgdRjg
qp5MUxkPjn4r7TT/Y/98xAz/8ih6BN1Zm9xgPUX9cxz4XF8MBH6jUEQwHbPqin1Z
3OMOik2UIXrzlSyDssyZOspC1eLHFhkeNnaGroYRxmEAqGrAgoObe3Vw6hjMwRKM
AIVqXbt0oZeu5z/09oNjFQH2RDVYeP93cbXikjOLBSg=
`protect END_PROTECTED
