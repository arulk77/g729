`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCkkuphnHf9c4sgFNu9YMH6CIAS5k9GgmgXH0piSgM6i
gcgt3zB4zNLDm/Iw4fR6/1X1zFojDKhQZTq4T7g6T3/O4NDA2rYcynNW16mYsP+L
VJ9LMOcGSZU9NniW+YQTL7e0QWwAiWQBVMRVfz4L4a5cuzKXMQ6KhKYi19xSk33+
KYgtx9i+SsGSE+Z+7Hk5oLlbUJ3FCMCydc8hRbeUSQygw2WHDHNRgECPw7z8cP6L
mRf8CJyrHpjsSzhqGz3E613ajK3lH2po6r+zE1ICUM4D7k0IUBnr/ytyChBA8EVp
4Roi8EHHoiGIYJHO0zHxbqD8hq7B5MPiWf/L6lmqSJ01Dc502Oga4zg/b8mzgEGg
t70GyCp2G6mX3lcvZ3IVGdfAO7Bvnof9SeyMPwPfCQh1OTi1GL7t6k+sCmQQ90p/
qNkiGhiRqKG4L0i1HhBgYnc/n/X9oieW6lj6dW4eA4zeOie9UK4KgrLMTSj5+Cc6
Xq8qT0oU+Pleo8vwR1KAbXClqoWMMKaRBPw+9pMus/1nElf9JQprkexuoow1v3kZ
`protect END_PROTECTED
