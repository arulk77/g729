`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1ae7tAShW9PR639DTE6obzV9MzdE6+dbmftxeHjKYRnKv
pDfsbeBuxvfZdAJ6WIYPEaDB23RxJME5GKGkfvu9XEkxKItdZjaF7Nlzg9g1SQkA
iX/sMrwTm7zLHNwfupQIXHfAjCG7/sq5hTCZuksdLUzMhM4LAWauEWewTtz8D4Bi
Xv+XJWQJiseRuQcW0YamgzK5/RLOmDfAR4B93sWrCG7iRF6G2dGQHN8NGzSbu00g
JwokbRVtTE3FerWTj7mGVzdu/rbj1mgskBEwBKEDUg43tqh2yhmx+KJ+bhQ3F+4W
bECoqsOgZu6hdZpDPVL/u2+mP6yra+3iJyhKFO5YGQxWVVh/zVNQg6XJ9UCx03u1
716C7v0Wa0W/FwrCXp5jtJlo0FnkjZXLZSxB0d4HiGrGuAdKgSjAahQRzX5ar/lH
t3xVrahOEvUUo7uRR4mzKN6gZuNFTZ/D0Nt+lv9gfNijwwHZ9o1YtBiGdSa5Qt0+
`protect END_PROTECTED
