`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9ni+f8tMjZi1DosUxlGJqVYZ5roKyPl3fEMnHRO4mP9bKYurdlLKhBcDTY90HGTS
1i3OmZnTUotiYXlM2VQ3dk19uANBfXBnwrhJfVrPqDuhjtC7dpYPWnWhKoNk97Jb
yVXHTqc5WAiU9cXZUX1+MCzkH27YZQKgVuC0zZF8qI1GgQPLbNuSCF5WgQwD4I0q
rWpttNULHUE5FTLtFWRPFW/mdFgiBrtdeQAby9Vk/ArYL5NpGdZyZBZsVt6lhV92
ipYKqFKtmbK32Bvwurdg2LVXHcVV7+Lugq89KZs10vKSxidOFFZxT8zu2W/WElEK
`protect END_PROTECTED
