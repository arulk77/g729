`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNQ8ArcaoCq8IzgXGZBd/5si834+DRl/uCcK7Wj+1PCI
CDFmCTYtdUy0mSRJSX/VPOGf9jlN13Pg2n89slVGDc6rNoWVg7+J1iMeyLhnHddV
DvgcTNeoCD/lZ8a0gJtCI3MKnTEeDzs/1+S1zErOo/Ehv7Yo2UmgUWI6XLaGkiK2
br00jUFe++ctuaqq+9PllMb5tBEkhAT2JN5hsctgA9YSs7ZCT4asiaNT56JutFvV
a6moZobL96dHnMYlmCjp7fOcIUpnie/IOKpbiE+enQPQtKYnUoLK/IP7JqMvv7Ln
tY/0GT8pDUFCx1L/I3bobceFD/i471ff08XFYKuaRugLvJb3HMOu01CEPWZatVbM
ueC+xgOJgGbXOaYMuHSxaMHlYRNlHRWOf0Ek8Fnd00nQb1IHqiMVxYhok4bLvd5T
qalCoOC/qtiFXmIDEDYwAHQUAo4RXnF1cY27UllT0ed/TuCjDP2TjQuwr11NyWkf
2FhLERMo54LGORVxQ3XMfK0tgzJYlNJDlaokIABZVEsLDxnU51Bi5F3NL+9el8tY
qmSdXbB2QOXKbxMKKxmZ64MKDHx6ZYMSJg/NOpXgGo++DxmlpLcpsSL6p5M057KJ
BwfGV0PVCbb68QWD/rnbMdeS30r2lCi9WvXJ/FjOIFXYf7hPQhPOjg1JIn2OxLKu
`protect END_PROTECTED
