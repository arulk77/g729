`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aa+sc0qsJTtuxjsKVD9UKUv3COSYONBaIrKo/xsHRBck
dg6Jd3XeiP+PWnFY09KCBOM2LOKteYFXGAcgGpLV0Wr0MKPJNPS9iLAfGOEpl5Da
DH0jS9+bvMiKgvjEV+Pe198L2I2QbGmZi7NSJdw3VGzZ9MtcZeX4a0sR9fW8hPrd
XEHOQ/2tx4yuCiOhFPeu3vpIijeRevl/+KJXvlnai29WcbktcKaiERoDTzEDYhLr
1FTa67sNjFatngj1O0afL5o3rlNhLnmIka/2l7aydQ9u0Ux5nKnNuwz+nwzDzZsc
La8HvuyGuH9hhFYeEkr44b7tjhQ1qt828IPxj5H3k8wLjIa4PXgKjJPAZ9fNU8ca
5C9ZV2nLxlMakjYDWVHOQ6tMhu+u9CVzZCtlMd5T0Owqo6WHNdB/1LofuhQjJqSC
YCJsTDOf21ngQx//V9EEyLPp/x7AlrA61agVJ5eQrgHnweB802QqUxMN2c57BbbN
EL9i70JFJKXe7X/GOeG8FA0XvGDTjUTS+NnD4fufgydQlHEpxvv7gDQjvM2oRJmx
z3/m3gcu9+kCtZHX1NpbxWhEW+euA5yvUwosfrp2+c3nlSSCdYGBicsZlc0fXV22
JYrxF0kuMiGLWmeffvbZuuJM2Cahake3/SOSDFkkONkLsKUGarvdsWArUiwb9Ahw
9wey223cnzg1qQ1KnGlP7SFch0BUpu5eli8GViHBoK6h+I/eTyXIrV69MkXgol1c
QgXpDcwBryP/66WGHkYoDH73kbNRDLcQY38wpXwEdcj2dgLtv5t+/Z2b1My+gfKv
NhBza9AT1Vx3Lgu2jEgSaxi7gK5anKj+P2UrGFkmDM0zVOeMp2INU/aROGi7qW02
KCkhz/mYyDmdGy4mSpB+4v2FxNcjjs/kMJ3MOkxptoXx2nRngP0mC9qEz5yOITfp
cz+272c+SJ0ERhz5Jy2iOLOWjcn7Ss9m8fJBobUUXoN1s6OthSPM5M695Gy7J7X7
MlVn5BzqrKKquHsq+oDqxxVRQYXEShVp1JrsJM0wkF2Kwvmm6NNOvB3iXcmc5v2d
UJe/xnCnOsC+Sm1ZfF8V9zktZgPE0X36HcREBAedDQu5+URkDSIz/q4JGx+RD05K
6oQWun4FlbaiKUfz5Jy3BlqPu1PNt99YYoZ1wPKjtS8iOkCaF1EH02TbtSOIQWE1
Dpwt/+ouuxgHJuTh1RY0rg==
`protect END_PROTECTED
