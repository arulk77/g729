`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48UiWhrwgEiMPOQtcnHgS+g5kCGfmxT2VIMje0qB8ECB
xDfbrfgyBz4gRPJe4w6JF5lOaI3o0Qt4arEVPwTOO6lRGdgvWBg6hTMzEyB65AqY
ko2YAsAedvA3oA3X/2VPKnURXkFuN16x+WY270f1TXRBxfuFWMc4e3QpJj8ggufq
lCApJf+PIoTIDkOyXD/AeFDAxN63wQt4e8qOQCgr2SvzHHR2TkkBSXm6l8epud8g
uKEXdFQi15RJOAhXSXicvMCOcZTfz+yd2Mr1wtEe4nxF5HBKhpoCTqwMGdpcueYK
mq6cECL5xucEL7F/ZWH4mJWUFrq0ellP09itCkAF9iAasUMS2Rj8Ke0Tyi8HbiHH
MdB2jM7H7Et64pmjyCBvvw==
`protect END_PROTECTED
