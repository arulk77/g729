`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SXE9K0VZdOMCcBnRIEH455UFECSFOCpsPvbhZwsfjr9O
NfjiAygYIJZZqKJj8rCezAtTAhnhQd5JynKhna8H+3T/5+F9RN7lXiEdQ9qbcDvV
N/4CQMvUnEhOTLm+qDn4c0F6Gl+Dyg1zgZKF82L3goT7YAVLW+74L6ZrIgMsCuH5
XNvl3FF9KlHM0odjRxTZ0PxomGDrLLlwN+Y4YzZdbLrU7I4T0p/pOTlGBUWLhzab
uIroxB/WL2+ZTeWBMfbpycmjb4abRAYDxPuLmCsYERKY0k2PGCglkr5LGuI3Qa7D
RiuNbU0/v689EXIziaAwbgknOXaRJuIAmW2uD9VZnWT0B5RaG1Plr4yu4O0n9MDp
sLq5M/vZtJf4T5uyVlo/Imh215hdNjfwjUu6DVkRGiDsyBj/QAalRJJ6nUehxRjn
y3zD3GLtiZgQSQcHNWg/p4pQ7EkTnHsKB7/9yGSVemm0BhhE4FfijC9fIT4vnG2K
Rb4D1HNF6PSVnX7D401yEvlCdqg/Fvh7rBqS1VACkeUzJ5HZpvkPwIOl04OzaOa2
pJ+2pj1JRDDlGD5YbQ0uM0dlDu4RfC0ADJIyYfsY51scF2taHE37iBqTpB47+csR
0PFzFEHDWbArH67jrBZ/NJ01GUY/LlAXslqdRXnnrWs89CKwSkE8K9VMtzx+94lH
NhCO1V4sACGIfyw3hwfmFwhMmRZ8pcHFAt/Shz/BOFr48RGIgHMk7w/VnWY/oLMu
UGLeqXKXmh0cq/suepw9fi32FC+24phNKQ3PKuv4uMWY+APMPCF47+sJc7PFsO7K
6YeiAyfrAvThPc2rAYshmCJRIE3h1L1YNkdjbX6zQc7bBFGzrQOvb4nSiOK6v04S
UBezTWvkroEu6ICTKYuCiRG8LqtucDEhpE1YbPSr1ChEnj3Zjk7X4UEXyOz0iZBf
bubBoBtzAgBXj6JoMWOAlOND4CbOOqp29C/bUriLig6moob8N2B4y2uw2/BZfH3k
PDlxIRz6VB6+L6A9VPYy3W88dInyax53h2f9JGx8M+2IFqGRCGEVanLw31CdMaMA
/rSRb7iNywea5l9fISKd1i15nqyrems2dgl9l0+OHa5aaS2vqmADDOeuYySQSQP2
fx9oxJwsAqHmcWLqqqk7REXpXG4hualtKPiB2xvI/Lt0F/O3UiKybrpgvvEfFqkp
20WcwhrjyxGvHdBL/6r4rUs68wL1fN+s20bsxkLotpXjahgGYv4n4FqwwFbOEoUN
pTGHodOFq2g2QwZvMO4fc2Sw4DR9PSQl5Uy9VM1qXKOV7sWubUjkGh8sxnaict6q
+Vn815iYvAqQIDIUCHAqjPqkPkEOr1tQbeEnXTpJw1AKq9srotwGEJJe27R1CTGm
WdIpbsbPxJE7lS8MRuALiWeQYtwi59nlILmQSE0oxjJeCiVfRF7PaUldlCDTq24d
lJ8WXvQTmXAFAI2A7ldCLEXyomUh9IqOfF5HEW99WF6H6O1TgJzvP1lWzezlLUek
TgLjqmjpIdKBK8c2xYFpXhKZsvUfuZZq2rg4O5N1jszSbtr7GV9R/Zc4mEfY00Oz
acuwHAmMJJWvRcpnJBdqcbMt+h9+XFwp8098d3JFEGHrlYYINZd8pnh1mA+JjWB5
dmPXwBVCFDZklYzHptKkQnP1ACaTqVJKJdUWlxHqd4O2nkAKGgzsuM6GZrkEMxpq
7s5ANuC3HJW7S7XPu+AN7ds4Da44BEm2WfYSpPxtakONblxnlGhfTLwHh2vvdLOa
FM51mrXn/qr/6/lkQzhJoYGOZIJq+LRGLZ+TBUmh2Xvtryh+J9VTwa/KgmV2nIho
W482WezuVcnPsMcH47D/NcBQKtrWb5X/7r+OLFbdJEBlaOhqjgCZhdVIdvprFuPm
wtnuL/DPWoi1RwiGbPhmMBnrw0MWa2vhPl/M9h8/A0wKAgPGLdDNGtbCJ9mTHLhD
JCUYi9zuFKyubbuEiOGyioPByu3kka1eHdnVQjP+YgTddRoDYy1PKIwwUtNUkai1
jjsV0+U3tnB2MpWEVT3+EYoz9C9FqCzFlq9Z3uT+SChyQUrgdNmpzGZMmX9Cxvvh
0gG3d7RTrJyg6CfYHls8wq6jHlGKCmiaTT9ROxU0LM1e/01PaayEi5PYOxOKa14U
Gy+Pf+n2p6puGEGqR94RbVJ2dIF0E1wlBnxXh8i//0+uEy+QhRWiOf1zHsn4CTsd
2SDe3jmEaEsQrNKJwic0gQmjtQqxqmmnQiSn+uWfbQGuACZhuRtnAo8Pdq1wI+VF
3Yp/03CP/HPKW9K2iQHdDyko54ZXlcHO9X9b6ruXAs/TrwLwjpJ5UuuQMWu0wKE9
me1n7CovJfeuh8dPc8/RSoKtg2UabO9q5sEditXkLbYdfUobMiMjzmiFdN9w8gv6
y5qs6sTqLQC83oS+eqXchqBlwaOIePpxsbIdkuGNngAhchk2wMvtGT9feTAapP9q
rgmyPjUUTQ+XIABQiCDuzP+buenKmZrtWbR+bXW5/mDnuk34Y/DnO7oFwuYraUhy
fxY96ApWbGjLxMelkBjTzE2luTTzpB1iQ6jmRB0E0K/h9dFc/VYdy7tFa52lnxER
pkOVTe0eOAYgfTlPDJqGTNCzZYOfuKyZzlXQ55Num93UJrcVgft3np8zcP3xkyVB
elG69P/QUEpZ1PACPNdES/hINiCkkNRbzkqqDjHXXu7YvN8OGvl3sWgYfsgn9Lik
tNwIm8kfS74L6pII3KbEi6erDsuRe+cPFbcXFiGAtNgqfi/8uCyh8z//EA7M5wVy
u+sHbCsI0i3aM2VUHMjOx4fcEzN3PUEVQBR/FxNcjhGlvcbyH+FtLTCyVW35R0l6
UQ8bXYvojMXaZ0zdCmWBfXn60hNM7Z7rrVQ6c9RznnB3eU0AOLs9m3XO7qt2ws5Y
2Z8SKZbsmPB3IENNWQhlVXSAF1H89ePNjiIQn+MAiIxYeZCjYtjNYhNYcS5h+6Cg
SkTvpbn9bnuMeIkTZ/2webmltK2rlXviNNtGXuQPLZrmAjjM9GUJGuRSOwnbPLW0
OeP3XDQwMtb20SZalJT0krDheph2DimUNxDUUDrkDKrxneNzmoKu2qysn7Hznlz6
/9loOMqBMNR0mph7ttTIrfoxC9Ya4iMte9MOK5XS7vvDJoXsYyZy7ppHXhipvouu
23fANg4mYiOtOJ6HKaC/SBEW4eeZOb/HXDt8DWTqUY9w3bYPAQVE245cDEV8xADH
l/aiBEcDQ0g1UKejb7uSn6Nag0wL96KlMnqGBG1zfuzL6jkoBA+j9TLRz3OvtmTk
Bjr7TTsgGvyeKKR6aoihYakRrGf4M6r6zCpx7rmt6XlUd/BiZ/bH//ZtVpbfj6Xc
QEcy9yUjOLfnbLB2zYJcN/Mz1CROWrYSLQRpoiafRaz8Balb7tZ4UjMpcos7Qaat
Xqcy7o7ECzjLef/PPDSCDuXytZo6FVTraNloZ0l+oxruoC7pinCWFo0Nqv2VgaxK
yztBNyQOySHAzTAM7aDefoJ8w6y/FdT7wZr1kpdRyoEtOZTWu5F2w0Y3jz2PU09e
d2SDSb0O7oM/JYtuQ4I+N2oNhkKthidc3tYeemd6B49Trn8TEIW1OYD16jfSp62D
oZ2feTzhYqgnCf77cDWJz3Lps7mc7x8IoahUAJ82wDl5HTVHZ3VN7eYRg6s7EsfV
zIqhhVtjH7XeEJQ4Ja5Gufo2cYfbDkF++49HFRmD4umfvgo4WYRP4fSnWLmkERHH
+E1M+wvzLT0AwSSreZfXGkhUvp5DpnlqlKo2HVyJgRzX4A/L/Z8kVlMM/gAi9rwZ
6RLe9bMIFHsZvREmMAfo5yda90YbpBmmR0ck4HCCAhW5vi7mLAakCH7km9d0XpTt
SMQxUK7p7QiSd+bEiPY7hvmDw1hhQ3ETbvfs+ekoZz1YJQfUNoURhvaJ+gZg3cUV
gHZhlbfrbNNLwsXXmR1GZjQtgZbylXvR2EU0InxXCmKPrCUGrwtZULvCwFmdBg6m
DoAsPFjL7drdmdZjOwgtFihiYccEw1NojDDl+ufIRJ4NVeXy5WllitUZfArg0DiL
C0vzwWEmXBmckvzK8E1Ww4anq5kmQYvqN7IIqklrYsQ=
`protect END_PROTECTED
