`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kvq54R5Zn/rnHOCQo+aKTAnekpb+Ibqzzd0EqTuUVGaRFQdTYt7KhPy9GACnOGS0
2tY0zyTfmMkUTEcUBcmhC2SnmsVOCRQ1kVCkKUdpuYUmyk4ChzgH4gpklstgqNhX
FHcjOSVKEWbceLzrlE7ldD60EI8b9FOFKZQnDrPQuZ9g2kgxhFgdGLBz0PeGBU9x
nOptjqhPiZd6duRSInUzEB3WV6hrgnFF6Ul5samb3BsQBLPNvVGSKZOhd13WPDV9
2057I+Fc4pqYsMZvVP4bSC6AaH8U/T1qgFLL7lVCOSKIwDJBsqCjOTqjma/9bx6A
qwZFJE7We/E1FMgDSvrNJzjuOQLgjWTwDIFBT+8bJfo=
`protect END_PROTECTED
