`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
c6NdHFqgI43tvzVFaMY4mfTaWwzeKUI9/M7NHyCq83RTnofpolP70OdTNmwpP1Jh
DWKyncZpF2p0t0dIHtRJtxDiGiZB7H11YysZ6tc2j9rQ9LXRgZE3GH/B02D7meU8
LxYsMECfD21wzwTLQkYiIsZbketyFvvylT0m430oNHDvxkV9n/HXrzMIShrpcZYG
wQuaM0Olo4GRILOLYP+TmXPlpOXSTeErtR2d7D0bDbZKaHyWPNvpDmfOYmbvqHvU
`protect END_PROTECTED
