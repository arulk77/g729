`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCn1rrEijM1S48zKWtqReuAGND57xY6fThQydc23J6Ti
8a1+icRo/moclgJ59oGfsTrfVDqzUN5gpnSrqotkRxMJXn3NznwOKcTi6XrbQ1eH
rxHSCJ0E5bTbq7wm3+42ixsgMY6qr9fFgfV5dzon3cONmoE15H2ABs9Z9bNsyxOv
BWVYx21/UuLv+XrFgJc/Pk5uo7/V9YPSx0ujgbN9crIxCA9m2Fym3F6ShTxuZ9cM
EohduTWVQn8xtWBKolerlYosyxFsHcHMVwuH10Qu+w8VfBbZEwhTRM4TuHDCAU9G
IBv+Y0O1b8a1chlJvwtRctLykHTw2tO0ezaqMNsUMMGOCxhwLW8IXhAYrj1hMjOw
FLMszR7Ba5e3nS1Ymm5zkVh3Kjx2X2Qu+WdB34S68s6NImn5yr4COpO4rb7TQWbJ
rch94JTazHNy3aN6dzxPxdNLa0NLyLmB4ZBiizxCz/U8DKGFTx28re7tS3Okk6Jp
`protect END_PROTECTED
