`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIswA+jfbiBb/uZ0S2uAxE7TgbVG0ob+zp7Bt92koq8M
vX2xWVrLUXttXORQjzMgt2dIaSRMkPaddZO7dWAeGNRv3C/pFGhItzlnnAG9srPV
6zyHao883zhxW4XgBNK0EU9WenbH/3o2zTfAJ22bJ6XEbQenCXXN71UYQ3b2r0Sd
jdRRTYcbhirCSOMjqyWpC4WtmwHg8nVf0f/yYzf/kl/FV3OTzwJsMqhxvoRHfKah
NTRKVPN+cMv6oANvArE8gjvj3SnfaJN59lx78NavAmRhMN4UNC/XckRxNeYZxIb4
9RaHPcfmRnioo4nkeBmGcizFbsOxiCgHQ/HXPXmZDfwX6J2Hs3LX+ErOfT6zG/TC
ATBDe/I56B0rEhNNkEKcXhvJ6YMjD1SlMmRRin7rhYitTNfZFBNvg/m/OHq8iLy9
c2XXb0Gxvv/o3YnyYe269ni1gcXhwTlNKoLYBmZ5S3+zODkIhCmXWQ2nG1NvqTJJ
/G3eNfdzaiBSoCOc/J4KqmxXgegdwWiZ6QzOnwMkC/wvBj4FDXC/VBBlF9ijHkO9
`protect END_PROTECTED
