`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNwUdBz+TVgh0sGCYOUtDt7LYGXRbvc1GkISsA96c3Cw
c6d+HyoyuaSaS60Bs6gdcejTGz448mewOhAl4foa31/2eamFa/mo+qRwpACubrXf
Pr+6WnOFAuTW0A1UGZSXlTDIbWEDSAwVI7cA2mcZEMrJtJOni8zJnmwupqKdykhP
qxDVveTYeZVFfDHMmj2v1o3lOI7koT1wjW7FsyU1Aa14pi6GBiijdt6L8B1XKE2q
`protect END_PROTECTED
