`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aYyERJKvLhHPPcyV/lWjJKsuUd8NPZuNGjeLFeG8wRYK
lRz5IdeySBVE5bJ0gd2ZOpb24LdKmS4v6LXhCPrR9KJd8ujn+ypqUrHssVX7eOhO
yJdinjjTW5KH90r5n+ruP/utUKIHJu3qs5yYcbfgX7LG81TLCcOW4zzqs+0qNskA
VEvcO09AKMUIRf57bw/VWJvmXPbUhkn1vJwE9SYaVkQ9FkfPrnxOFj1mqGnLi7AG
RLPS7rA7ZQ2iSUdQtT7Hb3bYocFkNyNMkg4QgCGqECTBufDhHpxcenahQA0t8yz6
/knaE8JmBnNxRd1lznOLkI97NjVoqEVpmER8RQ/FW1iY8H2h2eWYotevveDllMoH
qwICulwIGzY028YFr/DKKfhUAlebcStb1w5UqqGWKGpO/dLmbYcLifImehIL85uS
OadoKy8pJVefRvGHNg+Qy5M8kqbTUMuL8HtZWQx8uuIVufJO6rVwe3Goczkon18M
SCd5SelKzNGC/B6cApa5U6RgQOcIoqWm+KMH94dM7y/bSuotR29jVmGEilk5wGK0
8lTP7HNu6SNbpPjlQvtk3kFQR2ESJ84TWjLYkXyMncEH10+O4FzEqsq/Eu+4NDGJ
F9wqMKGlRZAg50nkYYNd9adxxm52hkJNbSlduxbNd2YWyDLWvacnZlompIDL4wad
V7rPSfWJxVIDDCzjApLzM7euH9HjTkMQ55VHkSx5opUU1sWD4Ait0jHXHeyQUeLN
t5gNgOiABRTeaBJ6PFZIkVMiYjVbS9SEdQsL6b9jLDVyzQNq0vnlhm+xXV6eQQgo
aVcCR0d1LDm1usY4Xy/bfnbRuqEEw4t/rbjdck9KlCgCLJuK6PE4WVo7xm2ciGRh
fGbY1QwGxU9jVPddh2vNR41DFYXTQY6k2cJxCC+6g50ivYqM/yUp6nRaJb0j/JOn
xSWAjEp2yqkWduRw1Ut/ZpC64uezuo7WfTWm2XTMm8yzpv/A87FeCi7CXPLTWC2G
9oUkNYvMbPG0DAfFWRBjhEN7oifijiZEasNr3hllHRvTd86NlP6lXOaxRF0xsj83
LS8pr6xlTke1fhxy13QxWysDgMibinmbADf+9U3h3EfP/+cBOiI/B/I1a61AqitI
DUA9klpSUmp6qOIExCqyZ10J/qpFCPOvVP8DoomM8gDtqFlFGuUu3p/9IlvCV1Ze
3x7IJR+8EW64ODix3ZuxCin7q5rGRnqI3KKaVTzi+goNCez3Tw6WrDG/BRjKsmAv
XCmXgvf+0ajWCsgMYTAoBP/t+10w+uTqs3GnnawS/3o8HcVjJ22km6Pq9dXsrcm2
zxrIb7NVjLrP3TfJyuZh8+Xy79hxIgq/JCvuU00JLNNlvEyrNM7Box/dc3atsXHN
2/umu8OgM9uPvOFWFzDWwPKvDAeM6c+akJXpCvB6d/B+F+2u//HxQCihU4ed7p8u
ZZuJdpk1iuKvsL1BxD20xOnyu+s4zbWePkRp6lx4waUSfNf3G/AaHlTl7A8IZlIs
sBhfMyHkmAK+LgsWGaQ4RcjDR6kOV+9bcrRnJcjz/Bk2La0qVUETJc3p7y+7106+
5R4rDSzkQPhvfnv9unxGeGLEl/1VpGebgGGwpFfxotvfRblTqktli3p0U4VjY6e/
4kOrN1d8MeMBMeWmdPLw9JMrcYMlbcI63Bo8m1tzrlwjr55EgISc/Vf7yugGaK2e
XsEELC0Hc5D5X45L+2JseNUlREQuX5eFuLzC6YBWDw4d43F1irKGhJBck//IHXGY
iUzbWlOhMGuxqV7Nd+yq4i8V+5xQ3kzW4X1uh3pNfP2vw4K/Hw5GdqvdivlfRUqr
QD3+2EqQ9yXQDwxIXmCMLw8Fn3uXIUNJJzJc7qGKPRNVjjsWugMghwqz4lvwMw1x
TNI/mdY92+1B+3HWAlBqcoUtx9F3TBHhKUkLoSF7t0k7t2Er7tWZciHKJJYEPNIM
XYiauVcQEDKy54KXHsK6j+WS8xz7wZwM4/hUZlnS3s3kBBNeDfsAWVDwAmqxZXd1
7glX4Gy2LWVvUERBAWcN/mqtr7ohAZFH8D/4HIvR1jU+F1ZCnkF8hhdboHmUxVZ4
yHRrSG5eqiQwIQwoTHF7ejtpFPHxJFPZMR24faDp7c0=
`protect END_PROTECTED
