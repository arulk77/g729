`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C/Htrp1EV/mZAWe0K9D26hHHjdiyu+LdR1t1riiKpwl3
i/DUy5EbdjlyZH92juI/z5eumTbHmvTZU1sPkru3VTvvhK6pStaGrTr0C3+5pnnJ
6lgU2JfE8PQK+jXyBV++uhoQR0nJXqaPaZ0h/E+mwgqhrDqi8HjQJ58Tzqqi8Und
SDsdIs5px//gTYRr2etSNLbZpWuZV5qeEmQckvse61EZ+B8y0DJ3C5ADJnFmulNC
RVNQdCzuFOv7t/6T6EGlk5qx+m7rnHEYGXP6HSeqdl2HYGmW/dR+mH1CkFY7h+oo
fmMl+xtPgnNHhsocWO45yYXIL1fQUApbkwoo8qlq0PqhBphp7VWUmUsdLocZM+bN
`protect END_PROTECTED
