`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/S3Z7S4ZZjqnnj1SeUr6tG4cunVhrvRWQreZlsk4Kjhq
wjKawjt37BTFd2RQj/GAc0PUu8W+BpFjwXfnIE2d8q44wOPVr0zVz0TvMXO0CF78
+Oq21DCjdHQvwPEFWBaEo0BowBHEzLowWPHPeTaaV9atPXOt3wC0nhI9NHPE9d6P
1AA5+LXb2E9e0FkJs/wcNB3JNLJqr6QC4J2VMPCE2JE+r6HnEYT/pMnhIlB1Hjgl
b6omhY2ho0swpVFg0cnUjRUzHSeMX2vxuE0y6xaP/Ou4gb70uxoWheW6y8X29GNW
L/icvDOhvJhJuwSbBeQwjW6XrItYD+/9VhN5RgFimFsoXGPcl7sNVzhMpPAdP7sj
`protect END_PROTECTED
