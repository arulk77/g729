`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMJqP7Rrc8Njfy9qQ28O1gKULXqxx/fQ1yAPgto/eeco
/dnLQFhNb8c+UCB3rut+HEdRjqXjpFQ1+mIMrJdluiypb1KAKFGZroRHPDx/0/GV
FuhhL5SRdr6o2Pl7zBHWI5gqredfsttLPR/beFwJe+0ulrVbd3OwKcm+esc0yzma
roP6rGmXT00y3ZUP/ThaVuLan8lc4m2CZVtp7+eH0u3E7ShmmVBJDZHsGYKbL38U
pCv7aLRMh2f/wACk76HuIAdZQXfK1sVGdjt3CKYosxjpv/4ysCgeag7g9Mr5IrLM
y/kR3htszpM+Kv4tkVYrRI2NpV+axbka01nUgVLkjQYmC2zCYVZL9o7By6h04vvC
usZk6AtaLvK/u/ADp1DoC3cGHp6I9/Be9oNuNSizWWqc2fl0HIK42Fs4z/mp3hwS
9MJvL3/kgCopt0JhVt9MGj3CTd6JnFDtbWcHsFNB0QRDCzxA7cEL894U0z8wuHhs
qFh55GPa/rg38og4nNPwEZDmLzPxDgdx1TkJQ14R+i5BEv5ia71lQjlZM6j/xymn
`protect END_PROTECTED
