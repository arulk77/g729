`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMcJy/7boUM3tFvBVJSiW52VKs91DOGoab13cHJe3Kg3
Jky838GezD6Cp81gthK9kDfm+dcAOnQuDXsq1aK/aIj6Egzr9HwZbkayxfcu6XqP
e6GlcKVBx+ok4frm7FML8/UOnXjKqRh03OmOIe4ddyopy4HBYmcNTwYKyX5qct+k
JAAPmm/CfjDFu/MPNXyfAHFcmcAOfJ1CQ+wock0jONHZBfHgf8XqM+rDjSL3E8cI
hvt8HSjj0BvIqypP48ocQWqoH2AOVBV5IHm4X8honMdTYh698vAgKB0UEb4pOMvd
bgRrwAWzFVLxrriLW8+sgzyiyg5IdiKhlXJ4nahluDv5j0bcpJQoh8us1YOkg7Bn
KlZS4V9p9179edg4zRJ9nl354D3DWMipZ7UN4HBwjyba+0Z9ou+APJazjcx1b1Wd
4Xu3Clt75qMBSh5rw5T5qmgBNfp07VxqTEwk8Reo7fVXw8zSsE+ynQZIASCqz6jA
we7FxTsXw57LDMT8PHqQsiN9IuX27o9FLZ4HwhispLhMSaRGUEkzGhAXFmnQyah7
WhheQtHtopG7tk+W6/thYtWl9p0ip/Cr1Hqho4L+0P5rOqkg0LaZK1t+vmJcGPii
uKlf8jJAWxL5YClvGf+vbwHoXOjpjciSzFrtAj3/OCNT5ULrD4oOOGH5pKEvSxUQ
`protect END_PROTECTED
