`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KRGHv0sFKGPL+twAf1PbuIIGYdJPRUBiP5PA3TdqQHsYT
AXa1rcIB8HXDb12lzr/5LcUvNyXezuObo3FboKyMsJVi09oUbVCixoDw69MxhEpi
H640LYcbZ53P2gQZrOGp4z9PE8zwZFXEFsxIdNvKPZfwetvnw/YYjgibd1HJBi++
`protect END_PROTECTED
