`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKnMW4r32PlytPnfBxVg3H7obSRrVLPBzjmUwXw3ISIm
w8gyIc7k8jm3RVZY1zN0pf+bFikic47jwhZ1e+TjAmKg6x7KkSeLLIj4xSs6rdSl
XvAwtdZpvJVIjIQSyqfCdiB6GPuxyGSHFDg9Y9ZaO9+Le/tjtZOD1nh/lReCQiXL
IHJ2rTWQ4j7jioObyrBRjvk6LOWOm0sL3URHUwzRiWziigPLSiLV53fwOcWahOFq
pnuRwxehwBAFV2ukH73qSLCAIpd64deSvuTO5TdOH3Wo7kkldYbSxMDhl1v4QdMJ
P+QprTNrtS6M72YWsMHDaCQKbN+hlkUKt5kkbjq0HD6EZMRIF7uLLE7V7koKiEE2
bu6xSF56FuXIPNrO5OSVk2bg31qNmZdbqgYyBbZ+pQJm8i1QjpZJGRv4SASWMUJy
xdah9/QMLPfFyw14/9e4XOsn2fpu5BEavxNsHTWfUFdRSUU+mg7wSIM3qFEOkxwr
mG73gZ7viws6aP3e4vPSR2cv71JyVDxjGIaovquaxT8b6Aw2NSyI1JsjC9uSJT94
`protect END_PROTECTED
