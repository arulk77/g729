`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C3/XYEf8FRRvFke+ftL80d8ydqnUjTOhjNurasd/KEsm
RF5ojm7W/9MsamH727KeE2Zer0p5w8/EvkaVlNB1gRcUZvpeem3lRvOkjMsaKF8a
zEoIA6E00SsLNOxyrIEIxfL6GociHygzYlXd9ANTNn2GmmQD3JOsCCFv7lU/J+14
m0L+as9Pq5RtVoF2h2ARZfG6E8K0w7ShTA9z3LoGt3ijURA4GvB9qTTC+D2LoccT
xUyIBQxIE0hAro01NAyT56rYoCI40rak3Sd1eL4lq2rtZXy7rMvwj447UU2EbM7x
tDh/OBSZD93PhvhfVKBlsk1JChWLRcIAsQxa7OiLkhPG+hC+VMH54RdS4uwdpr+U
BDuNTAJNWWpeX2tgQQnfWrecR3c3I8QrLIQhBxNLfS60UhZP0Eg4PPU78hGbvI9J
5ZNjhKX584fiLT9WvWCJwa8F+olfR2Oa3twyMOavDX9x87Niv2CLAFyxleHoOXel
cBZClqA9uCzDC+ObfsHeDBx6pd0n/CudnGbRArlq+oe905W0NX5/I+F6v1fH3m2b
jALNR+PM6md1ueQMRlmf8gFTzqJlPVT41uif/NDWBd3KT1Isg64ERLj7/jaBPS4r
toPuLG4dP2Mwrn6oc7nImbads3VyQ6LY/E4DrcZxFYGQgLD72mNkPUXKlUtsp4tm
zIUgU9DNkbACuum4+oRbkXXvnvhpnlsYbT/kCF+VTYffVE+PXAAsseviCQYuexPJ
jAGZXapO1mWlt0LrskjpLpwcH7MGib241oQvhxvl9lwvDp4jtRkxfVMdeJr9MG+y
2W41FdqDo7w5Rfk9NLV6LHnqvYXZoAspK/nmRoBJ598tYR0ybOgUll9gQx9GbXCB
Sqz0iHkX1AHkKjZTYOYps2sXtmCCwjivEJCa/Bkc9jzi15HLhHYmJIlJnqFoGZrE
Mrr3qImtrUqREYJiQxfPLulFr9JwfxYtBPWd56mnRMLKJF+RtkGGSIuRo1nIQOhq
z98Bpg3NMdduKXWdlpHDUufh4gooD2OYXKNz2KNmkHfSZh4L9T3tcm9qfK7ofrW3
w+wadYD3B6zyFZ+Pi+yM5m7FG40ycPvjIwMIZnG5rCXrbKibQP/58R1qT96XA12u
xVIHRhW0Az+VXTKUEWOx04rPY8hYGpUcRFvSeTzsBo/vP+RpVa5x5JRusDphnGsG
Pi0tc81QkiG+OU617Ldj3AwbvHpkfTXoziTR91sOYyDiJE2hPp/BItNzrfn5kcBG
SsLt7+GeNrsHTw7Kahyf058FqdqE9rh2RJZZLYSVXbX+9xLKJqSjBsMfjb2TTqag
uUSsodvCZ65K2OUf/9HDbaUmNO6eX+YXjeBS1S6Zc9Ri0BzutDiPWclq+ROXCKH1
rsgatQ2EwFRu/dSQN0n0fNl4HlxSwIrK26AFdyfOFtYyjjKjzNj72gLxCyws2uGQ
X4t/ZHF8Jpd6q61KS40mpZbqC8CigKnzBlM6/5f6UQeHbTnVwHJU8OKmV9YnbJy5
xKOoWx03E91xrMMd7rMdVEgteGBxpVEJPQnR4t1gjP5xo/eFbjeB37BsSORz2mxQ
2UCR4RcEIQmqDUKkBi/fD9v9os9iRyMDlgtTCd9nw83+zmaV5BjS6nI8mRaGMM3V
ezO/hopnovOaTqnIyiowFgPFRf375AP55sokK+s6YYAczaON0RiwTiGoEyLazwVJ
7RLyOHrQ9G/95AmRQLZFQMcp3pzaFJnrHY7YwdQD4y6ydWA+pJmRHQlHnx29YGh/
87TymnrCCUQTHb8/LOoSsrc5h1TKGHD++A9cGOaDEKKP7kkZei1b5m+7HKPcJoIh
nAqWgv4ZGOF4Fd4zLF5hz1rVp1yKqek5+UlMVjJHV/0a3lg0ZdutoqNtPHZ6SGii
qKDmkGgLd6VqXiDmCwzB6pLuUdkELi01JUAMX0EGiytVGedhJjsuAT8WU2wFss7h
Iq7UA8uokMv00U2EPRLvTsJ8fVvZfkrO9cpqYRVBwziR/WKZ15HIxZH0Z7Eqzi96
wEh7EPN+2mURAWitVZgxV88ucVbf+2sHxKcsQN58+CGfTG+4XEUnGPlp54YUwLaO
eLQxg87X873gIC3hkJM28d13EB5U2UfXeycVzu0NI8lmwX0z8uWJDVCvEsAPbBLS
z44ShRXwwt1MNI1Kb69RrWS7cBy2sqy0THTdt1E7RsFykEU26qhW+MSmH5+95Raf
yt3xj34gIe1ATQu6wp7q8wnjpE0FjPISI76y1bFUI7zDT38W9fb7s0c+twxo0S8Q
M9+Oi3td0pHk0GGDmM+tc0cb/HoD+1AhzlWPx37au4VHm5i7CPFRLGJnk4Ojc7ug
pH84fVGSJq1WvkKZW3COVyr0pkoSbQz1y9sz6YQt7oVQQSJvkR4i4rttO96zakXF
ll2pUfGfIuMeDrFkyjRkc7Dgk8LiHnYBNee/Q6Pmba4ZmEWkhg1sWMHcTk2+7+Ca
fQPfRL3MQzUKObdiShhjHaT74FsTJKWc1g2knbzpzjKO3EKGc4x4mj0xf3hR2e49
bSVfhW6KGyy+4yk6/svzsfXYxm0o/27DfuFGCUlO1Yd4avp2zIsHHpNx5ZZcYDyM
ysYq4dlsyWZkcW4G977R2ifW2E+9euoV+WIjP5DFGwK2ZbDb4hefFJHpiCZB0NCr
m/Jy/rOdP1xXT0kFI7f2vM1kLwIQQLiQc9VL9CQHzCvpdLULUcXEc6QeEtnS+gO0
wKrJ/mexnGJfk8bl5Klu1bxfnGzpKlnJwxlgQM7AAU3L/CAJEYWvnH5xBVmtQa1I
UE1vxfIT1uMYBszirIG/FDc3zepSU7GXvgfz9DYI1igjbQe1T0QmupYA7rYJykjr
PJqRg5JM9OJmj9vPKrzs6rN4eO32qWd6YW666OA/2f6a+FDwUpfMwQiG9wX87Tbz
CP0WT1AQBuT8YW1VypDJRVB3KNVljbzTayN5uovonfMG35wqcyTLq2NVC250/nbB
bCx8cMNpD4u2fIO2P3OjhDxS//RxYgpWpKpzOPA4v7PQ50rTXd9YL0BkCV4IcM4/
9hOZsc6yKOkNfAA8La9J4kDP/zMAMA/OboDJGVsikOamU0H2RVy8Y6pV5pSvDarE
nksLNhgqHcY5UNJFZEO8xsyHUAnwZGQ+KLp1o7w2JTsjhNwLEewvb5pO8/sCuyOw
5Ar90T/S9yoHLWEU2MV573lKQA9pRmf/i9mei0Wh3RH5zzxjzODueQWVt7c44xAI
ASDPU3W64CzS+vz0uy9uILtQqTVD1Gx/h6Z12CvHwrJsOUbLHHrbtV0q00lfL9+a
6Ma+rwi0sIrSkBlwYtbxKT2KwhJzW2Vf3a4uJPM/lQM0Fc1ayq3A3EoyQfYdf4dR
cfmhcHnsfRFc+0XicOXKNX+n9l20bdTN+SLNr+1+fWjFzREUBtgx8CXE0tiOe6jG
jynixcUVeM5H/HCovtj8VcF4aLiufpexBObLtOFdWfjIzjF0RlLE8Htu9bpMqte/
U0jgs8z1T6kB31EdU0gDGJ95Em2JSqdjJnp70ljq9YyqINPujbeA0ADAk0gtS1MY
UmQXdtgXGuD8oz6Lj8bAizm3G4LXHH81a/PVYDvW22psMD3/sRuGH7VVgkzD212N
SMqQZX48+P0R/6Q3hZyJr6KcTQDnnmcVz+igSaekph/shpRKAhKxFSE7P6YX574P
SwQJ2r9Pl9gfu0OejplScxiiFlyCJPRx7YCh/5IYy81gWG8Zmtxuw4n6qqdI2q0f
q9hWTD+q1KK8qadGrulRWXsXCVAwF9Vj15nrSA2DGA70flJzxaU+mLG+IyP38joR
UpDQIwbe0pZl3mp5EfOfD7gzz5DJ0iNmwh96GmRToEAQ146l3qhNzNtdFYxex81Q
Ud5KV6V30qGE6UKMVQRZxqOY32g6khWLOBreRlq21ek/LBjaSkgdwxt7E1jHvcQT
NTMPqTXqqx1f8eeoc+lpgTN6lGs3rGLydOSR6ZP8CfRro02sSLIJVk5QqCjmsAhi
E5dHOcBl96SMk8LZDK4L2vH8nYVWD003t5uD+yxQH5oRUNuFIw5acjuOWI7rw3xZ
AMDe5Rx7B2uL677CKrfdzjR+Mj+ygPMv876lp2fxHVzHMy5ZISOU4kj/n4yqcVB5
TioHYpQv97pTCxTmGiB18dxcOEqwnZoXUSZvAPUAJr4/JfcLHBAPTaOlDFGXTnxr
y+AB5Ca2clDs476Ycg3bYnCz4p3v29Gu1hAGmQzQbpS1kfPKmqN3lXYofCQh7j+c
sUW7997ZOuzA7dnsosgCuiUb9APplbJeoiLFSpcOP53JNaiD3h3AZqiNjJcNy0o4
S6IwkCk+WMvkcWdRXEPg07xOUJJZByyqaBK/wqv29sJoP8x3Vf1ztykDl+NCsr69
fihpv+FhUV6YV3N2I66N9s858TEr1tQfro4FXXW835hGuvyTFJTsR0SJlQ1ICyFv
LMagPYfkHCICPGyuSv/naWMNMUmoTu5qchH6QvQECvJfMliRT2NQ6QX+vrYUtLYL
ta/DdUT4XUFvLZmF+p1Jz/jQIDjGQ8JY/+rRymJl5AbzTJy+2trjwgjlp4GSamDB
+ZHnFySjgUaqlf75ArK420bPUzHLyD04rx0SeoPh+1Vv5Xa/2EAf3ZlUOq1RGsdl
Lf3xWHuQfC3sbuBMbFDGYBzpbjUXY/G+BrarCeA3gQbp1sdb56fIwZ7Fa3wdY5N4
+QwKRYZRC3ls1fAJxzJ/Xv6EpAEnprBVt1070C/zPIXXygZfJOitzoLqlTZRKs6C
PqJ0symxrAgom6PpnR7/TEB5PT9xFauobEgbtEYK/CUoZRtlbyI1/l7t5/Hoc2IQ
Q2QsJ1fG+0ENFJzIyyKX8r0yxnmkl0AGw2UnKfDp9SoDffcFDK2acSDhsclWH95m
jKwFO8edoIIpC9qjUBeqquXiJCmKauG49DPALQj10eD4HcobgeINyZiHjbayVGEO
eSC1OC1D3mWqcMTvhD50S4d7klL2B8rOHuIZ4+LyjRTlZLrz0j6RC0wGvPN+Xh27
LyDv6W0DtpZICnIUIL3qM+1zC+a0qTC6tzoq0jUNBuo6K6tB5Wt0jDE3YNlyNiZO
QIvKIVHcxsjAlOGRjbmyGlKLONcGMayDJ47B4WoipKkLp2ByjhkBHmT2JeAtyzeu
7+IlDiWlvMojn9fCZClt/I6Ic/hxBVWSL7Z3XLSi2hqDM4osMrGnKUv72rRycCzb
eLJdNfM9Hu4efI2U7zOq3q9K+G4Pb4vW4X2onnUbDY9p+nZqJtxsXgNK8GfGe/cL
JPdN2K/BKkKoiq8aZxNuEdhVN8cgQ5KxZFqd+Byq6oPYWyKDb9q6GCKWlLtTFl8X
tslvyDtkZlXMJ+th0jWCZtiylp/E/t+PH9sPz9tQQsjHqPrcgRsFA7XGaNMrJMlV
Ci7zMDwGyHAZXK/FhNBgi/eKlK0J4/+UmW9jCPxjlF2De+cqheeHa1FIF/oGo4aY
0n39Hqa0i87RSr/GHeJ0Z8ySENOleDQobl7GBG33DN6aZQIEiYqVxZplA0Rf9P12
53ZTFGPlLQr348nePAoZBGmVNj4vRSPcRcBfa95LpsCoIwKGn/61lIS0CmFDWnOy
gV8o7y3NDnu5zwHcLGdpTPv0mbIoavTq1NFwQX5rvpxlfFDftvRK3Q2KiACeZXS4
bCEfxOr5QZbOCM37OHTk6v5IRfYYZLpMh/017FEE+a0yCwIXAwNlXh+Aegnh8C/D
1s2cYnw7axOTyiVdeztSLbIOonAT6nUnJXZEcYTgI+BDteQfXUvO2hmv6e8YYxnE
RAKhL9nkOWvbvcmGW69b8Y0jdtrAXZ+waT41e9wu9bGmxSYCXBtqKNrn/KU7rqpj
Jun3ctWmEttddGAil4FzpfPszSUJxlkk1UiXsMU2IWz89ee70SuIlKQ4K8HyZ5zm
ufm9NRDwxNQQ8rOc8+fCupjhMEJrCqANmdyc0nlDRJbUpM0X8zOaK68J/cCUakZg
sAoegMxSdAMFWTw98E35hq/Iv+HX97wMJnRgoPlAB5WKIa3oww6Pu3z1FjzFsaBn
UrYzx5RcATe6g+P4B7OwcvsTEZOf13zKpzCBeYm9RCrhbGT3c6M/40O8hNijqbyr
SfjnFO/Zmg22qNy5UQvZq8sTwXbq2S7bZj53NrSG1x9DEiid7Wd+GkT5qySg0cjq
TZPY7bM97AmVcnBk7oo6Hv5GiOr5VaZ3JdF2Q14XmL0m6TnBDDLa9hu8v7FuxiYV
eATLh6XU/y21sDWj6VFejLVchvizARZSPTl626OBpNh95fMZH25kYn+/RHZInWRf
RXOWdvX3Fn+WmXpqC46bV5zVfosLbSIc+925rH+0yxHPIciKqRIm4/XTMv9Ea7S6
2bqWzY7I3L/o/63MmmWCLc3SAt17dGLEfIYm8p27fP7ATEGINm/FmrtjENpNNkUa
B59i9Z5aLQHl0KwsyKSTisfA+sVMZxTOEZuLTTpSxr2KQfbN8nZhmd8bNwHlOXFu
Leyp/S4nHWEGVeuwVzsPM0d1ziEJzkfDD+tcGuPJQlNYN2V3LmXQ+/JIZOxxhoVU
IK2RGIMsbjjunhw51lKUtFOv91SSpoV1LgKSZZqrUmoA+KsE6/hmOD/Z4gOf6Wa3
ujFSpvHrhVzkil5lkTAT7Kn2AGV/uWpZCMScOzl2YifZ4DlOeTgJKy3i0oIaAzFL
wl/6oiUVN1GbQz5FhpxALYFUgi/z2615h8qpzoakEAteNEMVdqPFd+X5dH1nDL4e
OjeQmnjeSv4emSF0foiWAc5n7Ht7ICHUiaQDMP+YRyJ3B6iinmt+nju2k1ZRiixP
i1CMq2d9ziH31bW0DgnSpklejAG0Rcm+CgirEYQ2cfYRBN9Mmjf4iIcW2U9mHQjN
WRKpdz7yXPoDaUNIWikIJ0Ldm9uFSSAiELZQWljGhbh43GxM5451clynNPOZCBTE
z19Ml2uNj+PwPi64lNcvjkfH9hraqtLnMPOLashvzyZvmM+Ci1XTJy8uX42ra/CT
LL4qbOJEi2+PfcNxBeYR5F/wLrxQdCeP8plBqobQS6UCbH+4IfcN+BrAZ0+wyrjL
AB2O/5cejbjNvifQoG2iU6mZ46szAhWZlXTtSYcPAMtXQMniDDxZYet4CJ7Aw53n
RYrN2dludP6T3GXDSN1FU+FAI6Bp+dbv0z46CZ+51+lS5dtUE+YJ+PKE3gjB43g0
eV/0Vp4OdH54HTq6fxoLuX2pc2QySGFaRMCAXi6LKXwgb8mqrKgAvxq98twz6iFu
QaG8yACFJXwwzWowaySoT5UvzbPKN0mMa8MLnh5H4f7wEHetkp++qzqxop6AUVyD
SCQsZOMZIgj+wmx5PH1HxmspLuwdaoUP3dAVQCgXfeRc+3Srvojo8dG6pAUDgKG2
XtK77mBJcGXAOCB4StFPMx6fIDXpBxdnnCUB3OTDdEFUvYGJQZKKyec3ZwuYyv9T
useq5oav5NSjK9BvcT8eZJ2mgTYsD3jOdvgG7zc816jY4lucYFfBTuG9YreGdCeX
rz7v7B+YDQwVhz1ovQRQRn9RruO9uSH+bi/Po/nnH12GyE67V4nki7EfVG1xsCic
p+QPG13DRLH/FfGyCPVqQqakAFqu57hoPUgB2Lx+NYdrYm0fmkDPQzvfn+N4btHL
S+sEWZV3UlonBONfTpSdBez0V4qqZ6ARm+AxvZ36fbZV7kOvuHylUekMIXYk72V0
VBzF+HInZyB5gW+wJ77Rrtu/fxvMdZxfJnHMehuL9zSwpLPXIvD8g7agYJUzVbPL
9URRFursoV54OIUswdVB0NuSCY6+hwNq9o5IV2eoZpaH0PiNpvet5qWOGpKgbUJT
6jNW4aBh4pEqEBJhZN7GzmxyeYyWIxir0YjgQqjxcv2PpKPxY5KTOKlsX6sInyBj
PEqudYCPBos5bVa0G4eHiJ07/Q/FvKlTJOsMFO0JnGHeYHDOt9bsZV+e5GywuK0d
7hoxkhv+4tEqY4n9g7OuSDEkCCnpuwQTA+pvs3ijYVF5PWVj7wvB34PEQdO2yl8r
wnTjjyYNu6c/0M/OMcnQqnQ8QvVibT2fzOPC13G3F7SvGHSeWz3FxGoZmbKzJ5JM
oCpJF5AtnabSgcGjLFc6ypT5t/F70piLksnrw1bb4XZap4gQm5TFu3qhOO8gute0
CMdYb709bOjJo3dU5KPYfU9thWdF6oeAGmuqKcZ9QACa17Qagrrv4lcXe/ei/zWn
/q6DWhVYbJj10jj1KR6fuh4/AImYaaUIEk8/biZY6Wip084LmEqx8W3lD+lcmIgM
HQdN+SZMZuP5m42/c3JDA3t1Yf5tNXz+SXYXUn1dZqjsNjz5jdlrH8TSelQoAJmB
ZCMmSerucQAW2tviS6Fej3Kq5gHlWZ8i6o7GkJzDD+2VmGRMy/rgHsfx8YsQ1Zo4
7FhwVmazQVP1XDQbh0zWrMjqlJ6H/2MsCKqrDkNb6CnI+wn1wwTT6zzycRLCr+1n
yqgNwEheUnbKmutbxopWKQkOLDfnBNlvCYPV7K5pcHM0r2C5SFlzeAwblbgvuoSl
RXvTrihKAR1s0eOWkQ7vq/n05YjJIDJauG/AFAisItZsHijZxy7LG34dqlo+5GIb
zBE2uOJvkvajS6OBrAmM5T2lCcD7Ec12QqCpc3qZFcr6W9LMpsrei9dJvwgazvnB
LoqvN+JoN2ccnygLm2nFPcMNzBB+/HjA4GIUKsqDSlFHm00jeHgIvj3cM/Z7WGH6
wgzDwE4/HvnJ3hhcTFuwAnrQt4OvGx+qSf7hVPZ0kr0/MN6wLDdND1wd9oLysLw5
wqDXpe62wOtPTHXARQ6dwdo0TsrsDrI+Gv5gBAAI0xQRGGp/M0e9iMUr+bw3tVVQ
hp86oAHmWQxq67AEyNwGiZLQS6FE0ipPAjeYXuRkPx9EFqKF24t5DtmqXaTUjFJS
VQRVt2Qa84XZfOnlLz6FDMqUb98Eyn4BpM3jHPpZi42Rs13aur2PkqS6xgaU056V
yKmCalxd1yw6sxwkmb5tHMzlnPMOqTCx+beLWKkxNZzYPUgYH2HTfguxHSPbDaps
ZcMRDp9hBBNZm8ZqWbpGDlN9CDeyJQSeDk6Bzpvv6w9BbAYU1AVqbq+zUKXRzkdF
4+khY2IPvi8JjSCAvk/CJFJc/Vc4K1KCH4819OZSY5g0qfdfhWEGAedJgNsnAG/E
wO6/dBMHUv2nya1cK8jl4Wi9MPIHc/zWmP4eEEm3ZgzZzGliKtrh4G3MrT16znr/
zgI5gFaVbIED4ao87+OyqaUUy3gW64YKFBcImoIhCnmGew0R372hQTR1RcdhYh+n
pb2vdHh6HO13kqrHAyyqMiL43YXeHpbrGnIWMQjC6nm1FM8wPPeNAX9tQhFR8mUy
y/fR7JrWmbxzhVdvNBHO8X1SxD1eP0omsQ7gYT/ccNF0CMlTOPgCIp1h2cNhdAPp
JtPEfNOpfiXjyqehpPp9Fh5X8hAB34EiC1VmTcVUG3Z1+6TYyNFK8kQrvslDmKfQ
a+Q2DB28oijqz/enBaJyG/67r1dRHrTQmanDUzyWRGEDG3Xk0CpnstilZpMXleME
LzldUPtBh36YCCBG101rcher41SKn77iXC7l/T3AitoSTZr2/8FkjdYhqzZigblg
Per+6yMUFE8EH4d97jqZSz0XsIVa7chb8eX/iSKcGfm/KzJrYvNLUPtL9LifuIaE
p1DPjXNi3v3NEoDwS0NkXM+kLiKfig4LXAH9BR18Av1gFhi/WJXLz8EF7dPZnqbx
aI2qSyhfijkoc6ASSUPcgZVOvDmF/G6mFJePod0n19Jpc/TOwOusDavtbuMNHgTj
kMg4/EfSZElcXoBqqKTdnGNJWUUgWSM/su3J1V1TzTM+TH330hEv4ednrbZoEFfl
/0qWUzHP/5jMVPFMJdkRp0H6gUr2LXp/OWeJOZnrVgoEGJyQf8xeCQnuoy/eCxz0
9y/nQ9F79unnkWMdeE5tTXlzJNhXaUq1moYqFFHvX1wmmpZI5hNlT+zMxz6R4WEO
GoD2F6WgnFstZciusU7u/npUym2UWk57otelq9i6rXllyuA2Ob6xzqGoOrB3qwA9
3ETfVkwsQoPXZGuBLrlc882+JnPbrfAzmS2fIJizgG+SqdAfoQ/T1HBSqcgivzV0
U4D0cE69MkcEvkygcImnc88mymP1o9SdyWq4dZpkxvLeZjXM+p2TuDwj3dO6yisQ
XHMNvz/rnKDCAj56CYaNbWT+0qsFQ7L4mK7B2zL86uPfBCF4DEeFu6YQO+L0Uh+B
wRnJPvhnMPVb4t2M20aiJhE2e/vHdanpRDn16+iWHaPI4aLu+vmkxIjyPEf7HG/w
MGFBTTd08NS5wMzmsgMDKOB2TfWY+btPZm9Iim5w5Ct/gtbV6MTDxcErWkATtWVN
A/HwPeXvdHq7PLK8IcAXaUUdFtaKRp5IUSJkjhBQxdvqkKyOuKLPZxMp8y6xbEa5
knORwZYfXQOgy0ZXo2q6y/tTOvupKE2z/CDA7C23Gv/Z0VkFBSQmf96rD5vj5xXi
s4kCA1PqIdJRetFqb4Oc4H/bb5oTC+kcqM+AegfHrLdY7MIGXKfnM0I/HeqnFWGW
b+BKD2QUEgNZYESlnMRK5tabifZoDvdZ834Pr9CB60iEfda2FMIf8XpzSKD+2Yfq
irm1axhP1E6nCY8g0DsDnuJ2azLEmEB8MuR/+858+k3h4oYUEkY6gmmUlfavi1R4
rmOlWVTEIzVuHvTkEeUc0h3weK9bjqAP0wk5r0uv4HiXbuCCZ2ouQlKyspTFxixZ
1+gHjUk0E3SEUxqyKXw8Ef6/qv4gxPI6op+yFeWJrAHi4dz4ZEbgicVT5q/y+id6
aohAUh2IQtPwSmW99t4wBMfZ0ftSREgtw4+NMGnmP7Y2BVNgsI8mWfb7W9gQ2qWj
tmGlyVeM2EQ7+mEeKjUciOfcyF1SItdCuqHgkeEY0wggGrpTP+qO00sHGTCFmnnf
7H8gnenOpRb5QAxSSIq5gILNGVa94jzWfLx2i8j3yTua0c0Zl55SWYTTFF0r+Zdi
8zaKpWR2xhpsLcKFcNbuqt49NmSTlUU/84tg6dxB4JE6DZTDmC0/e5u04XH5q1Lf
IcGY3ZlXQYD8HYRFv+6UTtg0Q0/YINkHHjheXtUfGFb++hq2SqHSZB5bYC+RlGOg
W9LFQqKkRTHIqA3Vd3Lpnk7QbxQKK6WP6/BNpKJ3knOHWpjjcgiKfR/DT/B6KrPG
Hxra6DTcEtbaHImJULxHsKUMDkvu0uzai5XgjMme4/oKV62QjdKq78ziJLmeveYf
eDWXetcw1+hoKRWiJ/SYP3+Wg3/4/skSrRwyIcdW8CqT459fh0B5K3eXLwMDdqzK
5LNhtyIS7lujcE3TW/nY0Xeu2vFeTfhOE/PvSwEWpEim0gX2bttg7iwSZu0SB2QG
EJLAzbcpKj1NXsISjlF4EF4aQS7grwzZg2V1qNYo4+z/ZzmDzd78dWlzWRKBV8Bs
80pU4lsCFBfKyy4CfDAJq0bPyDbcpqUnxuZ8R+b1gxYXWYU1v1BMjUecZHqYRSYV
9C0sl0j4Gui1USitlvXyzCsr8ArHramo/Z5fmxmQwlqBkpxNYaJL8QQ0bGrs5ack
ghNZVuXbnXqTi4CeYsO/uWOmP3ZjqoWh5LgtCcDv07Z20VdDyUwR9GQ1bJzw/3tK
W1rODXgExKx7vOJh8C/1o9mGw3Ruhblvw3hEBIiEf3GcRv8cXkrXodaSdlUKRX/v
0uRGihWKgb+fuegQ2piqEmk5Ab2DOiHbLr01XUMtpKftDL9ifBouAuIuhZf2Urry
L3VHZ5zKxe3YvuxmRZFPFtuPUIUgWTY4WsV+Nivj48h8dYMP9U/cWYcl1nIsawIz
yzmG7sMkrCsyWN+rwodk7O5RhG2niw18NKOOVe6G2ZJlPvY9NdvAeMgFh3ZhOHH1
nnbIgvbkYR0/IpfD5p7K5umcZyqR9dZAj5e21YQOZqjmGzHqAw1H+v/F1dDVVmQg
TtmB+OkloOAMnf//kpajcBRy0Aph/KXQM8xIz64lK2Iso0pXfxerrqx8oTlDU3xp
i50l+pufQdMyR9MqGh+uVkOxkVjvF3uWKFwiA9gjF4LlXmiATtFxzgmq71zHbeyI
bFJiJmTJhepkWbXWpRAriPqVE/lIpesfNRF6klF9M+sLbvCWrohqWgGyAxEI1IW6
4yVC8qXn/2TXpdgw2F/GNLb04UPpzCtrQz+rk5n7uUXe3XrYUteZJZVSCDx59tS2
768nfb767vrIZKsbOi5TFhvRETbwdSaZZEwRuT8trwXITv8ehnAgfqMWwJ2I5GMd
oWpCVH18Blzi4srmLa2OcIXHo+IsUbfvZgmVKirY6y/c7PXf4Kau2V0ZKOGg5syd
0KimspFZs0jHEy/pzQuG1R5/cP6eax3I8O8Z7s3L1h7BuK324pB7c+MY4893/kHj
56PlRadR1+5yAXcGVqbaL66kWjSDB+8kYasl40EHSnEKS6qAKENb1OxvQnVjKAZB
DeY6yStmuBIoScMtb9qSqkJkDyjaga49rx+f1vwbe3R53D4x0wPWr7i/Yq4Z0LHt
mRHNYEzr9Q7p44J6riPq8CtCfV8GBo42j6V3SZznLoHmHQw0Ab9/Mzo1Arwyhncz
/qr39HchheGfnDJbb76qADCubs4gP9KO+hsUJNJMqvOHFTYkVRscc725ixrrgP0i
vjCMj/on8EsTXGEO9hZ8M5nnM39TB1Xqzdg5rTYND2ibf/14wMpiBzy7ynCRtTz5
tOK8a4AJHcpEGMS2IrSqpLwaiNfD3nGBTtP+mLEKq26DeEFmAdryDskkh8PzmQdL
QTenb6CRlzRyQrSbg86J0L5kHXHOligI5UwQCE9yuEe+SEER3ikHqz4y29lHqR7q
roA3/sK4kl3ExoodeUeGifXmJ1OEJjUQaTn6fyfmpHItuuIYPg6pngVoIUxw9GJ7
f62G0ujLcpci2luuSlmYkgsRYQj8xypvWtkauwEhyB60XMawA175l3NfyTcCluDy
VCD2q9BJVjxDjRjybGCaO92lgCaDsqQFqGQoBEmOmN9O0PC83grjEHgtOEALoLCl
T38pmVojGJRda1AnUCTHp9Bt8b/qpHiXr5lA5ebqs3bdBUHbzXFxh0VF5HtF290g
Alc3oXc/lpuoCRYJXB3Vp7jyPJWxiSd54gHkAtflDTRhcTluNb9dCXTlMpgMTyKh
ls86ftdh/1AWpas1QgE3iVLIpFLL92QpDVsSbUDR2RoxQWP/RJge6iFfXNbWDlHX
Oi9YPT+IzFTMqgtZbJbh8rR3Utie4IGez4CCtMXaMiYXToWQV9mSObNM6Go/UZGo
Aw/DOtsmm62OPRSTTmFGnZCx0D4Lw+Q/RlV6XyaA5hDW3vOHsEb22J7f1sualStS
Z11Yz4hyssjbSEZ1cIwmAJbDtM7YDPdsgiD0CyHB9uBn3b4DhG8+0W0+XgltQexX
8+0IFu+5QvEdqMGLTlkGzHMt7SEzzjjsrlY5qj5+h6pzoE3oDBb6jyJxDtqlK/dj
55tyFhLmJDrtKKWPjuYinNIE7bVJaGfo7sS+Xot4dgdfMBQ+ftvxatEd6Q/PoEmq
0R9+8KWoSpwpiKxVq4SMxnW7chExkppQN3mspHlU+JtjuFAKLijD9KyCqbnds+3N
p0i6JgfThEz7qChqctcmy5SkNTn71O7/xZOJwHgE+Fpz9oHKOLbyQnsxhQwXwzRf
hGjZkviYHsgWQHgRdj4O4GnNoQgJISt2FCy1XlNCIJJb+hSDCe25H3nUZZvn2NPX
NHc91/5jnB1apSRGQJotbDyXrzjN8qiJUKwI2dmcpSzM7TmpzQItnb+L7z5GvZsk
CBpUBO2Rwz7jMBuy7O/P5OR8eXjxL9vGx20nMnJZY0evTNjp8vieHoiJDQyv22sw
9trxhID5EUatciGnydtIlNnVhP7Npyi3aVDi+vhlfE0ajeE/56RbEiEvfP2zz6+L
Cz/+mZfSwsSKREYlmn6FMDakssojpUZ7/6iy54qE+1NNtAD90WSOb9P4W7S7GvuP
z3MTeRvOab7YGKGCVbj/G0LKWrQxE2H/UpGV3XcryDPhx5PlL3mNM10l0Q5LfXD9
Gq6hJcgcoySMDzhRYIBwe6xejuiz+BIJGsdFMBTrZZLnbesivqLBYpM1HEVVe8TB
8lpGh0v9yMSCmTzRD6qy3dfPRqVPQJ51cUUMSnqXH72Tg1EPFKKwS4fq9KSaS0sF
RIIXeZ0KGGODUYdUmb0GdfJWX4+2a/1Dz44g0ri+YXaXO4YjWHWGEIiA4K0uQ93S
2lgOCvULbv3JE1rQzWnb8BK5Ajee0XvOmGUNfAlu8ri+bVf6oes/I7wQ922Ha+5M
Svwj4H5CQo4+I9IBI5r7Lh6qiu5RtLHMaBXibSoxyvUYQ90poBe7udA5xL//hyh9
pHTFUW5a3rkYQFqwHGkqJFjh7pWKYrX53LTfii+ZZ1xK0Y2GcALGAZ1fEFOyhs1E
9adfVz7dr5Ft2av0Wy+fwuUEmtlhDSYitRd/5VCRl61mKHXppmPgNv9BvsjlBsLA
mbrPf53iJ2yiCdCpsMdHA9plDeqz/cXl+tJ2BlgPNt2IvCbnMikbzwrYdIMNNT5V
x2NdMAyt9wKNiihGcleltwMGoBd7FBitcy+fVOMnBV1eovHk25uTWuj2KOE5Ygcy
QgbEwbeGRZlvm3/DOmZv01V6ApoRrkI7RESoJAhrCIUDGmsgf2njGxrhd+mCRYev
T0rS7YHT1iiiqay7wGXq/+nlhl0OF8Z4/ErVLzgzdUM/tcFFXujUiE9BUu+ly1/n
bV25hpstejMRn5zB84Debqgp5oftuvWandGJL1M3IhhBV11emcRqLoB4lBkWWlH/
NBfQGuTvAaGQjQTYtxSc3N56nkhB4iLMb3VCya0I4PlkDP5kPnNXNN4QM4fTDyx4
4WniGtnATK+i0nuOqQZ8a1uG2uYH/63EVdTm0Keni+Hc/qlcKmLWmTM+5jnAIEmQ
F1JcpOf4MRKhgEenuOmaIv9Sqa5jlOh503LLBpuiQIDmDiKWI3jKAIMNpO2uBktV
ciYnt72IDmic/Sg36t+ctakTNmEhuywZVd0wc6o0s9XKQLKWq7CNoisOAKA14/4u
BPASXa3oyONR44cRIAab1hhGRfqnoYkphV7EplQwDoMfhyMLOl7qTqdImlaOjM5z
H2wTtAw43xnchNcTl5acpEijbQlY8dWfxS4skE/U3UeGPNbp7pvGZtDE9uCjA3xs
PdCd64Bk5ttqTCIp38dsAN42lsLxKU1OiLWK6VtJ3h9gnAV36FwPiKaLEnHciQ0Y
9/Xh89juIsRu58GkmnLHN04lTT7VlmNaenXnCq4CJigFGKrYhrlCVSONG17VuhgO
MAO815xLR8Oypl3UbL4r3Q2O8Um/HPy1uRfbx4OK+QWewBP5bBPxC3L/pz2Orusz
XClQ8VtBsfseL14TFAHO89lW865ilaNiUSllllSpYxoHHh/A0uIJJDu4fTqSjdC+
RGu/8E6sUzU5nieIGHVP5D2dMb+gAvTyPIskU+76OvjV4d8g8U91i7K2dCbdOPsv
apakpdUjsKLEdyp+vOZOStXD21Gyc7hR8TlbqUChhpfnH+aqKqE61BLnH0TLJCWp
x4rZHYb4UcTRuGOg1TpGqZudSultu4FZJYJYRaHlJ9N7RuLfbUTUZOQOXlw9oFES
MKeWKimgvW8MKQXp/yFqmqZDc4FTFVctytng5RhutVfQdmA918Il2gtATfd2yL2R
mxH9NRYOGPp1IBFpsXwhzBBFaTA1v0I5e+kdhQshHAt7iecpeCXqO1HS211Y5yD9
ieNZWi8SMPW4Q0YR6RqaevL2UvaxwAUo55mObZxQj/90Ht8JmiSPoLy+dUbZCZTV
s7XtNPx615Zj2TKr0gOoN09wqnKfKxt72psYuE2GY+MlKYL7wS3S3YRohL93BgfT
3pp1U8m2bc4KzU5d7i1iTc/REzIYZQVejcHXMnpoPHk3RRB6MbNCMi5SJYaFALiX
go33NqK8VAzjchtRmnkrv5zLM/g3fT0wRvkRGal+7ujKlmwC1j3RNbM4RDc04g/q
tUiiPbOgq+Ek2JZwP5QY9M67szeXzkQGlsx70egYhWGgfRc7lFbH0B/VrrMBeZ4t
cSE79BWJIYVM5qxaH1lQsvgVrX2xy3nuBqqwX/aoFPn4owa6HXAVjwfOdsBORSjf
HJVtm9vMplZjvKRKqwdNUh0OwKPtPoccIEpAfFCPqKv7BZuHUJouEqElotjgUJcW
U44v6YhFWo9qLIwf273oQbuH3u2quV0fnYMPjikUR0vk/FhTlWhgRnel5ouHmrLU
CoCyl/HaXM2E/OH5mK+9yip5PBDD1useNUwjhSQoedJcxUZx4kmTDwJzw/xLnrhU
v+dgGb8b2QU9UAukPuLlFlizzxlvyP9wAbzEyWtbXrPlBl7RCF8aBdglrZv9I7ma
Aj4gLgjfnnJwsPybQxwLJi9UksCC9PfswSK/BVMip4s3fFswGbovpAF8Z0RE+7Am
m5K6Qou4Lw0LHjrsQEcTxVkcCNkJqXlgqON4brgE4AVTjtUgqVLtNGxIhXYlM3h7
ttGMDKtlGBR+9JbD7ACU1k6gnQK4luPYK0L/DY2uuINWxDH/xBiibJVqNbfLkrbK
/P1HUu6grZzr9kRGH52BX4SZWRCbs3T2uCrXw0CBY50RRpHUY503H5+EsS69JjnY
fiW2WZTyTkAOcCGFkqhgPTaRMHIAKf1K3NX2mHs3Bm4Guoo4IbTGad34/SljGDsL
OmCgou90pJGt/daNo5eTQ056TZiv94BJ+6I18P7plQrZT4XmA7n3JQdoahk5WB3U
ltFozYqF8fyKTwc7gTtuQdHCZGCw8Vh9LrIcXthre2AZtDL6m2H6WJACJhx2qNga
yVU7jrD+0s+Tzn6qlVPzRSujmasX4G7gOqrijcvOjwJlm+E91XYAc8r5jr3E4ws1
rKcchR+Hj8UWSn311sQ9ycv9zDY0Z+uvA9g3wQ4L7+uIdPdbpR7AvyYa6WuGOJ4t
6932cTTBbE8B2LlnkLoRCGBvqDge/vBL272DCsCin7nsnGCBo1vE0go+789pugOJ
OeIrFXHCASPwtdVq5/6F8nr4Or4ZF12OhJw1izwCROaTgD04G2sJXLqMYyHfWdo/
vdbHBieOdm2nrIY4+sBt9Zjd7Su9MMv+fQ2VBfjEhNIH37iI56yBZFvWyPigDO71
C/t77hKrfBZ4G9l23PF2wONaSTcOhhUKXfm+pw0JVxWRYlMb8eaeG3/RlxYyTiU4
EK6EGVshbojDkNnmN3GlFxveG9IOmbgqWZ+jNShExlOUhn0C/FfVx9d4DdmW1RIg
fcpr8bUTJh705a6rsGinYDweH8pTJ+G7yzCNSP8hBuUopjaX4Z4x/YNgYINXVCSF
OEa7tpWcQoiRlWHUyefD+Azfvb6n+eEASd2KbuN7UtkBKYoUStPyEpZDtQauC13f
VJ/FeJHLRYlhU+3DKCPo1tvXJoE5PBlpnZYwSfn/Chgl5IllrlQ2HoCI/X5GCEXs
D3qbMNy7vH7b0CxkiGfDfSkL5ukjLM6Wo7aRCHPdTqooP7CpDlxy5QFHQrmuUFWD
zym7LKT1i10tkwBEAFrA0QUVgokbKLa+xDlzb8wm5/CW/QPaKX9R2wEOJhYwfE05
kQ+B+0A226jsqb0WL6WweEBVhntVKRa87e27/WiQTprOOFpMdcLdHCJCsVUZ5J5V
WA48u+AkI+avlKH6jRGTaLCwxkQWHYRELF5RTcsrNb9DbbuD/d701ZAzKTYwURKf
CNd5gSC+mRUBjnrvATRqZbCLLhRMAzRlH312HH9BVn6/zYAmNi7HyBQXSZNGDKWP
WvnZ8bMB4QZhr7488pkPpwMxW+rExwNBtiJMu3Fb0cp4zyIbtSgO8PsJ8LgZuUkl
BUwm9fE7YTrarq0kOZG3Md6sGKBX7QMaLyg1NQ18OjUwJxXdp8O9nRNZoyD7DFPX
uEQyJXUt7nmQZh1e5zWthY/AE/oswWB+LHKmQafB4szKsOvmbkkTv0LWvORq8XMC
9SdcA9LKXh3uvWJv4hG6XEDhD1nHLX1OP1XTeB9Lnbj9KL31/hW9ek6AvaV5khX+
yb4vyzwhZYSt2GjmySxydNOyikVU0VooRbnbEeR/ggyoIatRta1G1kDbKcat++vd
FluLed+0lnJxh/NEo2BnWPJmtcZyklasSaEYLwdFLoK8sEZE/1TF0Jf+f9t+icS8
63xKj7v/gyHlALwCUmJqBSlkUlFs3reHvcYnS0gPn7KZX1m9CjOiS2tmpe3Pwph4
qeL8u2on6jez7oVyhLBX4UaazF0ioYGr0ShoeFSJmNrM6SL0oAj+8N2qTJkWj9Hh
yQXkIBs2tuN9s/sa+JQlRIe1Gf2MTfBLE7jPqXKGYDzGKC+XIDoLXOZDqJMg11NJ
CnRBL4fe8BfKceoyPCoeiIy+Efy1AarkdetKeqbLSguFt9025gQPHO4GlhzzVXtc
Kipt2QtdG/XgpnLvoF/PIAXPOi43MowrhARRTL7dNi/Vbvx0hh2qGZGt7m9PncgH
/UmEyccj9p6qGhXhVe1TQFW16rXqOWgx3FHHSEN9wlpNU6pLP9Le0UkxcS2zchCU
1QY8jrySwPPRSGKauDzYWEi/B83YzQ7eRnKr50YZvF/ZvSLbRFCAFAwqjoattZJx
ElFSp0QocMY2y62zWZXR852JpTNOCUwENrp7hRYma5PX1bf0/LSBX/kzxF+lvUL7
SttEo90Y9mfGr9C9X87WVobBrWuw4NWHK9n7Bh/yHIYfC1ojma5WeJW/2LFmHC0b
K/evkWbG2Yd9kKnUWIygNnOxmMCua7s8Ze985fTh4lp9PFBroYH+eb7BJEp8m35P
5avPdbXy7Z0/yCB5ETPrUSHNvUFKeMp/boBVL8bhcGW2DQZ1OcGKWHVgntny3coX
f3zcrO0z3Tyl1aSSOQiizqWlQGs2EaRgHOHKLVnqhTtscACjOOodjuJPz/inwc0O
fUQniZ1ccFTiDj5oNXBh00qHdyrTjM38euGzWNagiWV6Hx4srHQ5bFFvPs75QXLT
WdpT7wdAVo38xG6Lxdj5lc9xLuGxThBLGiTY6/nFO3LMFY8wbK8BzcQEZHmH4kUJ
WKGyGOg8G0czOMjKIEoru/3WZ1ja6b55FITZE4zWJVXtJO7GlSExB12nSvxPcPMr
Kwm+sxy/xxbtc2eDzqBaq3Ms0+1mgvzEWmvPhZeTd2xRo96CFPx6sT+EfZZ7Vypq
BK6WbAyR6wgjJ7LY78X53MS5WTtSKCgRs3BTeQ4EIq+GVBbbAtIcXdWvJYDlaRq3
t/YxPGrZN+b+a1BUyWneD0SlhsVXef2aZDAE0o4q5XbuPhQQG76Cq0v7fohbHg1w
aA+7jQT+QLhv2DnXlNl4CUln1NEYVxaRRclTrTVZqSmkg8qCUNrMP62aTZ5AQO/p
IV3DERD+s+ri2hXj6bg2Qa+MjrnvwyGXqD23nSeol1McIiTuCRofvFZSU7kdc8dl
2wssfdJJQx4RiWNNy+Ja4wJqDZB9fUQDRl3Mw+k23jcy0Ya8ByctChfO1Gm1OppC
QmVAXMfjDK/W7Mk1JykYkjV93RxgY4DoiSeGof98yjsAa9hOdB46E5zxUWPro20s
Z0/kLfDG9+5A1+Rwb9rQpa5AL3jLw2A4iN+yoFlnfn4ls+7/OAwPwu3FCJk20jqV
ljFzq+ZQngrC3/nMOdy6MpvnyEoWjXyps6YEbG1KXpV5+0xthvD6X9S81E9PveDg
TqSffe0oNqBeiG9rGi1CMIjgI87ZJmpWTt2ZRzzPep2glkpfMr0NxM0ow7aSsuer
l8Pt3Qw0VdiaJvo7h+gOsEpIjz6Gx3j1yEaH+kz5rB9zhbb2IH95i4sQIft3soPr
fMipYUOfWczGtPvn/fLOSts1FgTULmdd0124B6w9Cxbj0bzkgHSSwhl0AdHB9GFk
5auBsi/yxxgiNBKfiCU2qjQeF6wKNYUlLVrRi+Pw1P6T581Kiy+5R6zCpx/rvkgP
3w0VVr2Jd4yMNvVIIURcmf975wjKKF9eIw+DNy0jWQr38bgeL8qw7HW/Emr+y8BO
jCEYdhgoNdVwbEup3Ht23sDOUmGr06xy/CIa+Be0hsrKNxYcDg7T02KUh4I+4j1o
pOfwU8JOA+s8Yih8TFMSUceYLqODEPKQ1oLtF0dC41Cz9gilEQ+lEe7PvO2v1gBv
DnX0LXRlyIOtr6/AQEWNFPC3XlhcKE7sNVzAwy2V4yM4XuekkoXmnNROeeKLEJkw
VxM7//vhYlIVULm71phBETgG8s9osjX8GXPuVXeSdQ8AirmvWiUiT1Bc3qFgfTIJ
DZwX1Wp02GALaV0El3KyHKMlTkDc0Uc2TMrw5YIn+2Sf9k6v2+6sMthMXzbHZAGV
6/ReXy47iggTL/IrhdF57D+vTe6s8BGa2jxZX0hCBYDWrFlFuqBwIjC70Uqvt9H0
nQQgQYL9JZzh2SA3z0AjpwzGIPgmohH6fOHig3oOHb0elDoa8RqcVoavzWNowC6N
mi4NFeyfEDEtRAePnOTcINZDliNxuJG5o/2/GC5RykMxCFoyLiJzzQxRyrvHc4IJ
sJlj8N8ovPULdMBdEd/ti1xp6twJKhkzQMtmZKG+KEgJJMxjVCmzflxCKe40idFi
GLNA1m7Au2iWARzMztcLp6+n4WKte+WS8oaPq3YIe/s7He37nw5yOolFa+vyUjQM
UTRQk7qerqvts4vysRIJOrtbZa+M87m9RG59u4o1q/5LbFB1P3kTW4jAUDM2sJ7K
aNiRWh2fV3r0xE4ZWfQapy1dXXCAYjwnCkaK7Gbv/KUuxWA7Fv+DoZkbcom/3PyE
rRWqvcBB3f+iTCVDAOaGVEEajrKs2o5xb3jUuH6oagwZrbG+V6ep0yHk9R/VT3MG
pPo+lVErORmow/r03a5jkviUHY8K16MJKzmXLoFOlBQx+O4mA4yIG+VFwyYctqz0
LYf95eDUY8mOJaww9mOHxQ24N9VMxegVikHoqJcRjt9eCRmfnsPsRjZr/g/btSCK
qLHc1jYfqubRmolmiyiLErIzszMmBMZerYftU50Fcm/5BHfrhxSUkgf/deuRUZdS
a5VVsOdtJt9F6DFCSgjfOC3UdPVETnhA8Z+LuXH+FAvZElvkZq4F3Er/La+02SlT
pbDtkuZLRPvdwYhAZnw6YpavVQKVD21XGty7T7nk+2PbMGykNqzBdD9puMxTf/7Z
/BYF/rlo+IC+BnNfE8Ldh7utskxA8KXfa90jkutgA3MpzGeXBTPlQ44cFooLw4y5
6CwwlaAtf6HlAVGA4po1fLtzYNlUBf7mm9udIf/Xxtkr9VL1jP1CIRKPAzDxQpTu
9kUq6eH9c3ttecT19ow+bwwRNEAYPFEdtU0ANo10ZvvZGJ5Oe3OV8tMWw/oB2cIL
l3kTAQmDGVZgYGE4gTo4aQ/L4vcnDWQ0Ckn00qflArfABk+KX43xRGm+rzbicOUh
jcbFDwBaJYbkZbiTYsuyeJg78Sp3h+Y615JLZWISz1kKQCRQ6MIgbS+BuXLRYbYk
KTbUbTrAHRaD6fZnSpVtNu5/hXqjSBxBDnRDe1UaQ1iX8O0S6mcqAfd3SGzIW+cc
dNrFKtVT/J7faQQdBGii5EcN6XDeN/ycICgw0OlgsVXmMkq7YsOeWLAcg0FpQyq8
D2Az517mWXkTzouqrFrrEAbQs0LJj6jDt+S0qGiDJ7073Jr27eP4+Xy/CIDDQMPz
gtOhy5GRJ5WVYdPw4yDfQ5EsZYztjnHm5fvyT/l0JbR0GWE89hZOTWcswAqbcH1M
34PBUrgpWe91Qx7kf6NwV4bI71bWkmUDHTd0d4Ts91RJKnHtAvRhbEvmhlS1LEle
CE8aBqdEsU2El1T9KfwnhwI8wS3drwZrV+HSaUrGA4D+Q3ZwsgcmbWcFkki1JZzK
+HcihngQxPmvkGoXOr2VZqUIp7H/wobdjuXyy2O+6qSVR76o2v6+sB+Q5cOrA8Hn
krU3LDW6qLZNMWyCne6I4om3A53XfyYNF4fAGSo0nxSYeFEqRFb04Dcj7IP49cV8
4v7/kchy00mQJgiOb5B07B3sxt5nyfsYGQB8wGBEMyNQPUogQuCrEqPMBHXXRZ1c
Z+QXi5zIJ39pR+9DVHMPRa7vnyutfc0XW3FGGxzY9ZyRnL2nvuzzdaX0nqi2juxD
iSBTNRfKTuPcoPRfWdX1GcFlsoo3yOdR0+AFzodbrbMtMOz0hsfkEKrW1+/RELIQ
9j1kEDDTb/XPQ4+z01Nq6BhQB0dzBFnbfNt9GfBW2mCEC+8E93IlnIqf19lWX9dJ
M4sT8e6INHDeULePUcFnfA6UQwz5AHEMp7tDf+bzG5aQ9AaUt7/b3YoZZ2jScw7s
zHuNrvm/YwopgnD9faMXVjhuqAsBY4IHJKRwFzZZVNIk6fItdhqRJ8H+HpBds805
dOYhhmfYaMSPn3JiUX1KJ5Ld1weX6t4u+AEkMbOvk0+U2Xjcg03Qlx0yvBf9tmQ/
o04xnnzyjPHGlRfVyE/PFDqQMD0RkYnDTK6KxTpm9klnLMbwd4w15EtIqv5sY5wo
1gsKwX4QhAddCoC9wYhUeicu2OaVchuAxHlsMKBFTiyq6rggaDpCW0FfKhYWFiRd
OK0h46bY5J0jEk3VKuLvZM9K+pBKjg9I+BR95GTcZQ8MbieULMlszb+YK2VNuyR6
SfacJ5p6tzRxHLAoN1KUIEJ4oSXBBtgH5/MuAca+B/L0NXtA2zFIE/+7K0LuFhXp
yeZimaSQFZU7l3mcYyCaebr71Xk5ENsWviRTA6rPepFgB45be6wOpEfoP1Jpxlnj
8pm0SQ2KqLagSd6s/rkWQKPVUtsMWZ2apij8kGjsDcSJ2zVBft3XXF0/UBawZD9G
x4HLMgsrntNxox8K9fSsLFHGzqAIVuxFa+2ZdApRus8teL5eJOdXhzLixrK2l2ss
j04e0uTm3HOsGiQWqY/ixfJE3ZY4WEimQbypbSd7uBdln71ybGPdGAHlrBmrlDvy
b9z9KNw1IAUuasGovvdUzwYmxDcjHnu5l08xZ9kDPOVGDRgRRdvzlQLhSixVeqIA
khsln2MXV/SiHmuUT547x/hK6QyCWxXVtGqdxe3Umzg/pMVp7LhaEh8vjPp+CjPa
uZXPCgJqAQpplShbIm8fou92F9y5bkqu+3t8a0eMSkh49bOa0ZyaH7QoP1XSEYqq
OWyeIJXbjFhsgHttBoNx9UmteLRAHFG8uAmdB7AGFEto5RqoSw8XPh4fD7lost5L
YcguQxJfjZM+P5KKWkILAxFKA2cYohN+YkxdzrD4drSxGKEMcixVFOE6FjvCeTyo
SrznXJSOK8K7zk1nei44tiqzi9E1ghry3Qnw0tKvO1qqxXZDcnH5ZQhlkUgZYEvu
VWvca4H2kBEsGqSyqWhRyd8txZbv1KuBDRdVQQQPan5tZN7VqShVJj8v4e6CI3Tu
nJGpcxisnE+b441tay8/ZKTv7Upy5BnQDr5URPbGRY3srh538DSp+t61dP7C1CjH
WvsEHCxHh3JHLHoZdPhYVDwicHjd79XQxV5d9cQbcd2loCXvy/pdvvtiqOdOcQXB
e3RkzWwl04ZYsKlwWMj5lwPkXKZkQ4WPbSt2CGHCg26nsbctdLaZoKkc6TVZODVb
6QPOqUW5AzofpRrtarAd2bIzj0/2Bb510Zmmb0X5Pl8jbaNKeHf3bQVTWImcI4om
wgyok8wWVMqllzpfZC2f/aOZxjLDKnAXl0edSaHp8wA5guT6vO+WqLYBkhORYQhY
+pv/IpB51cPe778ShGl5x+CGRoF0GM/otQVaUoUs/QkIWVQp80pE6QDd8jcSqE0W
APZb1d4gOkhqdwGhvW7NIhx+IymIKJnR5M2eDK2CExKUDYGqMFTh1+slrHxUV4Yk
RnAWGnKbmnDebWdGTjYAHBQ0KDlVwfL1eBvym0xhmrkI605INEtGx8Pff2q7730a
Vp14OW3/q6TZK5NMd77jtByTI6/sGmR+B8UzjDXA64jiu5TDuaI+kwtOzOONAdTq
UggKjak15sEkRwIZI9baiY+b1qsxUEamp85paHel8UCcGPVv8VIlRb5H/x/X8KU7
e19Z1N/A8skjeuHWwnM38uh289AIYyPFXmwytq35mZzyZD4gp2LVUAGpzQ56dsIu
R1kBOn1JQLuhd6p8SBY6d7nFMqMgxw8y7H7ptfyDMwZ+ZO7IGx6CLAR1+FgIWhG6
BD+J/p6gwFqVdbmJ7s0wL+NpdyB7hqe3o49rBOSaoXEFkXvRxguN9ghfJL7KkH5T
0acN2FjP/iqtnTHTshaOncBjRr6fZ1JLvlUNDA3dVr4imYgpF9Km8JRmZDUftEF1
Hkf7/V8W8Q+BL/QSw+NfqSV2673YF88yEG3vOs+kuT/myyYf0LctQxem6DmLAc3Z
S5EGI0Ynu7j5t23YVG9aXrvBDdlxzG5jITxh6Wa1A9WWACQINoE5bxJIoh4dmi0z
5Vr2FLW1UGEABIOH7oE4JZX1Hy6eKh93viq3xWxaOHVmEOnsT4zIbIRr6wxa4pxz
ezNyMb9u1CbyD9cIH0pHXUMUlq8uInRrj1M8nItS5htjzD43gsNLlrcXrx9/J8eh
ZGLQwDyGzhBeLZZguOn2xRKc2JQoXotPxUShzzjOPsyWuHgUg328NlJucU+tHONA
tGTY1TkrXZXmyoQ8+Z95Z79mc4fl0SoYN3wpgaTJlyDNBV7v3o8ecjvifR3lF4PJ
ZzYQUgBgZsjauEyqKFLH1veO63Op5lfbECpyYHnxmF0788jpsWQyWsd5pWvagjoU
JovXV34HsIDvPZe0piUekemrFcoONoCYTW2UnSQRgJMCM90iX5cKsexTaHydS2x2
fL7kxukp2W85IKnuyh38g5mqFAfWEFOhOgB1NW8lwKgcop3qeqZhVTmcuYoV0Qi+
8KljM67yUisv/GPIl1Woaly7jEzOnHLsABo0Vs3ogblHZ5gES/mp4VOugsZNkt8X
TSi09hXCWv2qIruw7X1iwkBHNErENzUSk8HyLPAKWD8EzhvrQ3l3eI5ovYKtn+x0
g2Nzf9um0np4SeOAfxAMii1GmEHMZoZnPsXE1+J+bopHJ47O1p+tauaGllq+64QC
/xTghbFoytS1YHSoYgRPNncwutiOEcOs5Ts876tm/B04Ejn4Cv3VDBA4FxxQ2gmR
2xkKXfolCynxpErjzyVIF1TKfJdPxGXaHxMIZmBn/HkN2FO8Sk5lkKtlotH17t1P
EQJKO3RodWTUkv7WuafmLmpM+oMF/SKbvRClIzzOc7EvnI8qUWt40beoNWbEMQJV
N5+RjbnwyJNLVUjCx63U9Hbe2tsjn6XGwJeOtgxEgdUxp2iUDO8ZdJhdgg4sJvU9
jOO5Un5OyhCqVjgORrB/cNXm2ronsCXDhrjZfAvrojdAUc7sAXp2Se9kyBjRXRYl
rQbU7uF7aN0evIzIe0kzBQ4nyKU7yu15GH8XRbrqZRqcvK3jnrhzQkGEurxUvkzu
WtYIU2Ex0aLVcP5zpjNlvldS1VSLkXHok4CpKl4eCNcr8ACOmLaC0wJAu9mcJBl1
UNSeAnQbpb/jKPKlIWDSYDMmSk85GenNHIeyzKuR49e8gAH7mXoaFHMwe6hiy/jZ
9KHUtZyaUHDYG0xc2zaEFOK5jKH3Kf3E5PuhNWj2mhU/L91fIV3uunuziRZW9cKE
JXCOFTF2Yz+po32qJyG/ik84F79zPqoxink3/3zcFsf17AHLye5SS1V5wXHiVlij
xrSh0o+O1bwXKhGNCYjKwV08mn2uqObUAgPCtdRNw8o9x76mai+5iKSqYMNc6s+3
nxiT7vbHYoQhQ4xIHZdRbUdDVvBN34MXObNLRRnDEsqJNtyN9dC3dkzs8fPCq2jh
pRbwGUOPhfuLpErGTJ7yrIXMdKhJPGnu+N1uzVaOhPT31yV0h2HNi9bDyQ1XozAT
PsZ4KgpVNk5vU46RpoGj1S7nwbuttmzWBBcPseUKfoZSaUovzmHwjRxbpPBOvVgF
/Vj34bl7klqr+IJSnmbsRjBN2Ryirjx3ccKntLbDl5sT1zPCJiLgvTnPAA0Q7dBC
XUZ/hrFmxpA088tjiUKISua0RIzYqpr3VQCErFgAVXIUgaBqfkjPcSvnPafGDU1/
iXD6FLVnBkgqPl9C8MMOxrSiOPaRo/QDCLmSaqN9i4Nl6ebI/cb2wL6FLF4FA+4S
CTHLxvZUGmED9MRA8W4cXlEQ5Kg/bQHRHrT/67oBN+NvkWoPuCuwhcRv2butNk+E
aE9fa2vZ6+TuAjj5pZ8f1adoJXbnLwOv73bi7HEMjLbtQTI2bqg4tPCTqTsLxs5A
Rgs+0ZTynPDU0DxMDKi8mYaMPamQgKr49ClSW35W/GIxLvpXZ1eunXQJ5PmE0oXY
QaWdetB87B8H5D93kxiwTxf2RuBNFzsOdwU3KKP6oIiPTZ5SAnJGm97kUZaXiLNA
0Q3jQgQ3Em7/JnCVHNcbbFmGmZYQ3RunsvWDrKY0x2mYacXunp3fu0z1nZk3LWrJ
wTpJJ9A0x0mp+YAVaCODjnODWTpX9AH3bUOqoFjf3ssgH4mt9vFSeaoaSWJ5sNqH
l1mvbbAh2rIaVDbclJNgzvq3VvVm2qbpGWH6vHdCgxeiTnDkHYRW/08qimvSZawX
SXRtnzT4f9tvz6aAiFUKARVda6HcXbvSe+/UzbEEWAq1GtHVaSyubcT2LGiXinZ1
8Q/q97lXiTOfA+V924aYD38SeQh3VCSK1Jpl++pTdSxBxj66M1yFEUR2dNl/YExf
UJtkz1gmzeo1ar2oVe5up+1uknfCVonKvMair485exlaEM/4djUAk+3w+qYUujkZ
1j9jeC6v0Pere9qF3+jZyQfX50tRdciG9w9E8L2xAvam+eGO4SgpTv8V3KU2DVi3
rhCHyKIHBzTn77lyjAnidTpI0XyoLYjokG3csgeyxC4P6blVVMb6cHCFry6XRZwc
4KW7cZQ8wF/OoyujVWMpsqZIpdIqWRwxCFb9G/ycUvz7TM63v1ZKEjooO3qf4yNw
+tzPhebGy72aq3RliLGE5RgGrE/OfD8NsQ4XefqMHFsZCfSwpbEkVUW5m9b2lH2+
glzP1XBu8tyG8FIo+ILUjTJUTFKMxb1wgp+QHwaSl1lqkAB4aLj8/AUfWi2NAEIY
+d2tn5twHD3mwvjGKWywUfe3kD98SZHGxz3xoxi/ywj++tRYlazlEt9fsJCKTJfT
iJXadsKnVAHrssdRYPnwKLYZd+nAoqSrSDtX6ON0uRcMqEsU2n341rh+UNGcn7Lb
VQJFcr7hQOGEmBNvHGGeZ6pwZT48Y9JALw5PglrqsdDSEPXbtNL7iwj02Git9oEq
Qqx2T4pal4esOGY9oC1UbuPnWcrOJGZR9jhtN9dyroh9Wj8FalGPyZhbZ62ki4HR
WM1XatPHA8Bw3PisJkqSL/WEVBBUPNnO0tMEG5UZ31RQWivhJkTMAnmQ9CXBuQ9z
6roczGzHV3VlwWmDaVoHh4bD4U3mjdmYthreHVYK1AIE/G1vk6uPg754CcriTcD1
kCqeQhFsGuBtjUvP9MS4E7O3isjWpba3sZRCqkax6kb7dT1wOmjXoHXkqs5itstK
O/NaxfhqvSJtv9T6Y9mkSMgzXqRR8gzzJOgimxj5OtERq3UVzqTKNfsLu4yj3SjU
vBXS0yqP03EZtt9+YqrZhg3M8GNBSFrqul757PJp7FycVaOs/Sm76Hhgx9350GWK
KsaAZ+zVqxojDM03qX6+gHjFN5EtVvctQx0+/j5iT/CTQzPaYyVWS/9aLqS0j31E
Qm16Eqq3WmCiwpg1/IJNnokiZ45rjzXKUVvnn1QuQ+w5Emifomf9TZFNcCVqX9U6
RF0pM0E53nPKY3JijsMA637SrNUhSZFxXR+pviDClAF4fianZvgYRLt30yh+dE7/
PTgzZiGi+I3pg6dNn/rX4fazZUmWHHKKMARGQd4LSCSsah9a/jTAqpjxolDUxQUP
gGVYyKyEijJuYqpmluUIoC+ifa39XrBgLO2WotDQyEaM4TttulqIzUCtjsLVXons
7zRhB8Al5izV1OsK0e8JqcB9AhuPCEl/p/6+mpgMFcBYKg4JQI3z1BKKeo0bgvRV
SAb1Tv08zDdOqMZFtgmClL3MA3fr3gD+GfTxEVDMtJt8p6L+h+CARY3vZIWA8bpu
gj7mcNKWmHyHlVZvUy8SsA+nVuo4Ckmo1DNFvtl7VmhSSNftYAaZnmlv4XgmN9Co
mS00I4+2tIElLc70YU51XA==
`protect END_PROTECTED
