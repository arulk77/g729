`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLWR+5d6lfovSsGhxVzuRGlgdTKChUFtsirlIbhr1PUf4
429Z8uZRQhQc7+xs+IQuTjU5gDFkb00Xd1BrvBpZKcYGJuE1Fin4RF3uSLwQmN7S
g9SS587GmsxLpAde1AnejIZ1si6UUWd2BJ0xun+VKXQWcKEcHDRKCFZX6G4RLWjJ
axVM6roRcLVJuWUdzIE9qY4QBT0tZ4aH/lbcxsC4MKZ8p5re7G2tZKbMjmE24x9n
lt0fp1txXXfuBEOhUlljlMeCGb3vi7jWijq/iJjTIyc55N9m7C5gTPiTFE6lncln
ssy5fvurNTYFGTnt6vObVJU16aqrro7fH1pygb+X5nagWyAUTEjmSUxkeOvQrZuU
`protect END_PROTECTED
