`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNJjWLCDFoDyEgWE4qUMJdi6judCS1XYhhKkMGeEpuwJ
0fRu+xl0NIjRmC/e0Mo9jqxDWFFAvmOBX2nC3IIkMbPaKKaYQpV5Mi0Gk9aS02xQ
f6obZg/iZaQYCUtt/RPjaYgPr5cn4hn3CBfW/Ed3SvOCN02MxTLs2Qbvqt/0TCGH
eA+Vl+1Hin2gqIFSqpyh9A==
`protect END_PROTECTED
