`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NICyr+HJbUNce2iBTaXrennYCQqeTtuPQ+uykWWEOLduflC3x3fgsmRIrkKA2/Av
zeyfMn8dQsvZF5LuAU+e6Ih1BTZvnSgXNxqFRhmZPe7cqt84v9RRU1IBpjI4BshC
ADbfSWUZTzv1TeFslMHKLTxcUTK/JK9WwqWTDQ1L/FU=
`protect END_PROTECTED
