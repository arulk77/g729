`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6Idlm7p5xknE2zCJhJGFDJP0t5eHC/dHXbUE3zPfMxcPCCiSXmCM+XU0RJNTu0Gp
zi4S+pN/WSUcYVTiBdss4B6TK7S7kEk8cgASR+6QoCZbioTjZkf3IxSPGu7EtHUT
YurHRIPpQj8Ux4hkWrKb1C4g8i3MWEtTy3gTyop2XpxGs9Bw3xqApAku61VTwiiZ
6aI59Abd1gwU1AZpu50VpMbj27ge6mfAXtZJnI+IWQiGOCdVfVZ2yhO7s1uv0Buy
ahvB9I8HsDvmGqCrFVkFIppsEa+MK9MYfXCVFuimP+Kpae1j5Bzm9cK0IThsrtE4
AQr9ExwDTQyCgeCyW9dSakHcyV46wHawgyVS2dRWk4w=
`protect END_PROTECTED
