`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK8x8WIYWuStGLHon9WxRb5LhPZOJIWxIdHQY3feZjlt
OjikrjxlrmDY35/wUaaI0CjY3CYQtSR7DPFdE7otaqxht7/2YM8+Vyds2oxYkh3O
DUnVFpAibUIiZFY4792FgFjTSkP2PRIPgr9EaK9yzMMwxzXnUmnf46kJv5zIydpf
+p7sZHKQzClNFhoNNFEFz+HTROfqsJ7Vb00TMri4a9sUSTCdBXgoUDtqr8vNbsg/
WAQyymlHfWM6rLOqeezPR9asU3p03hkqSSh2aKzsusEPncL43y36A6lVfm7O575J
DzpcB9JsKaqdzbJJMAtZkKNj73VsrwXEe3ozuZN5xTmdszmCqyM5l7AqXD3vFzDs
m5gaF2+bM4p8iZbRu2ZGMg==
`protect END_PROTECTED
