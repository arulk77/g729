`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAczhxcyc+qG8DIb2wVVy31iECqLXapXeHQkryBLDqFys
kv+ZiHFO45LMuOU66iGttg10nRjPMjj1EX0O2KsUGglybgdTF0pG8kdj+VXSutL5
W4KOdlE/LLGJKQlDvxT0W5iE2/CHDHdaF8zDB4rNyEK6sEVJTqFJZTuF36z0pEx8
Hia2r5HrtzBugH68MlMN/kMbkhbTK/M7GSAbnt3MAkgGFFB7g5v4uJ+exbZtNncO
jY2KUJZbHRunbswLxTqxNZuio/Ul8TcoljU1oZIMhW7/dQOQPI14jDTxqNSnVFVd
gImVuW3t4ziFk8/pxJMQXBZGdAJN+HOG1MePoPfFJLKBZLeE6WiNkCtkBQZJwDwV
j9LIvvRSF4RbpC7VjHZCMlkMiZPL8vj8FwrU4BuHiqhx54Refm9lg4wsX2QBXioe
denzNhtBEj6G1z+BEV12M/u5KK5CwiiPOkeWDVjbYxKOG62GIvO8SDM9nou9t2AP
NvU0X03O1R33pe8LeVVXB2KgSDX0YqxR0O9lNO96wmbMOHhAebkxmSh0SC6efEb+
/XuTwzEFUzqBf1pKbSXCSk82HDYqUzhiI1IL3wtW3RSWFy8O61lznQaOQPmtkI1+
Qy2izSgHmQBR2KsIvKuRjeRO4/kWvAXFUsP/bmEH9KS54VBqlu5X+qN/ar2t5IDO
UUXoOSz5BtuQY7X7SkROJb+81UxVsc2u4RQP655/JNERVEXk+g2P8LeJ1nSIso2E
fiQlc/LSUvftGQ4yGV/1Ymze3frHoDQAgypS4CniOkU81lbM1TmVWYep9tIPRL+Y
l7LupCExls5btKrIJa5pY7eNLbdmJo3JTj5OsEW/2RWK5a9CR2eV6Jlq/24Rc5Wm
16XSLwXu/RvuYI95fu194yJSJvrFG3U2OsyY9uIqJTp+wsfnuygp6Ew8m6/M02aq
7jSWoqqg4Uz1SWBhHXzK3w4U+Ik3ui+4ClR2VLaFkPDHs4QQh1ncVwtLFgZuqbo/
fvWTaKNgMAm8JN1wnjDlEqAor5TPlOrTkJKWYcZt17PUl337LHbk1Kw8awuWR6Tp
SQUj/PDdDvh+ubOsQAmXDjItjccZx/PfRSg1BJXd0VcF6L2NfjHSPHyz79kLhLZC
zxwgT/bBTEwmwz13oMdwa87NPvlARzlNmxAEGGOqvulQ9WzoMfcc9GImFTE1poK5
NnMe3LmIbsmb52LsWVtHsEUwDK7PxeQ37gaf7pcJAXlnTKLy/Xo4t0g3OnZC7ECy
Hg7t9+TqHHfzVLt+kFr1BG7Y9d3F+Da1/moAMz9cJnqnegideqN5MNCeTQ+8dFCy
3ak6JIasKeTzWiJxcu57bBmSmRNzuJMqyciJretBpdUHj9RGguNKyc9Ht6kD28Ed
5nLh0q4VFJhjuVqtg2fsBPd/adNQTIwHH/pPlHziaSdLdF8Nh+5ShTGpVQO4h1vY
CQBTHUFcTyyDcDRCPutDGufVAEDh6s+jx3+Z0nDnhqqKsDW4ItH8LXdX3+zs2CkE
SibPJ/1k8xZMRbnsoybuy7sBzMpQAzdWjSkGi5Z8qbQ24eqQwKXx3W48lzXGKZcL
eYrOT9OMYY1YVMvPkZax/wBYWs4NsyIYajcJNvCSjFJu7+b5cyDH8K7Zph+6f37i
WVGbXsIs+Tbg+TwA6WNEHaPncSFB7mqbbT6EiP9Iym5X2EETnn8McK/9hOJ1o3ur
/vWN0Lpdd984ZyxFsYiVT4g3fBFPyjaNdPKDerwTx6cUOyg5j4voKbx5yuzsVuw/
+tirCqcqLLen/RHLBz1HqxSEqpvaSRUhKep3Wzpy00nCHGOofFdKO1lwNJxIZTUy
SWTozXUb+1OGhNp0KlsBXWYK2McmYsR7QOmWXHH3GDVMtXlqkecrK+w6FGubM1Uh
lW3iNMqHXTWxkMsHjquaLPsAmpMKUkR4W/hsUsKuSNB0+Qcn1pqw/uzJDFP9wHQd
eLXTpL7b9HV3aYEge2wqW3n+UdBDqrRSJn37DU4q9db5SgSrkxaGJknsTkmrLIDG
e/jUK6goLXLXiWZs//pB0CxCr6b14b/5HOHC5ilYPAXwXTeh6KwU3NqpQ6R1PCUU
/DVaxxymwu0Hm+Cg+sjVHisEa24sgBWhuiDyEuMdlJVCQNuna0/rjs43WtlMYKKk
8AyhBnAZQtuMjmzUW4D4J9MQXYcIziqVFihhe8DA2O98olMO+lvDHaNUJB8LXky7
6bVxw6TAnWHlmdq7tqzyCJgYOjXfzPZTXWAulq9RgxFv6w4/Ndq2oBAJbNQedfzQ
GZ2NwxFMpfKTS5RrdOtc69BcCgTjzd567RWUZ15uKrGFztZJj3UksIDExdtttlBL
ZOcCYjBRw5NXcN2o8lC4npDTvhgbSPnUUqQatFCQ+9jDGwQPXb050pnNPXWg8c/K
wX1lN0PYrCr+wnEfSgw6alvg9r3o6Xk/3QJsp6ZlyHu5oBWr4RHlxo5L9D6+f6YF
hwZtk6iElE7ykb/lAUGDDJS47q6S49GqKOMxuAtqAi4FoKObwXTdV9YT8x50BAw1
chykM5T6JsOvHjhq+sShAZeUjtd7svCsgTPYsMZ8Q/wvM4QRZ1E+/sOEmlaq5R4X
4jZ66SpyGxKwfoEqOH96DorUWoiiuKfy2p35Y8U1Ufb4NDrA3k3519zFRcB9KsAO
DJZeOpgQA9i5nVFjsDPRIljYr3HQyWJ+1VdQE7qcN8a5zDuka4JyL2UtfyH7SQ3D
JlBRRs7haqO8yPlM8ovAx4bl6Y8n1hwopDiQsRQ2HKOL1V965ioxkBx5PAPSNKCS
2cIaEDXcrNQ1DuIDvf7TsJiCEjBHRRHi9H/uCPoFwmOgPEhdiMK0IGCNGcYniOX9
yEN0DYZL5rnM3oscYVdaPH6UX0G8+HHM3qOIuZgx5YI4QAfcgO/62yFZSOCnPE2h
Ai0XY1BH+/4at4vhZxwV4JpE0VDzXE+9Cjj0U6GX8HxyhlmrCiBEVU5G69tAONnt
7XGuQ4msOOrubExPcUyeFTeVcvZOdvyp8lRLgO+YFfnJaf43W13m+fQdp5b4MYJj
PYWlyWNKGM3iA/kAXWCBe2WpqBqxFJ/Dxulo1iDgzoExMHnjTEvhHMKdrABZzlaM
bZz6IFeedo2Xb/BZ4Xp7hgIcE4Vmalaxp/QuUkxwJbWLKVyu399GJrtaSpUSou75
liKeBh7ZRQNPZRHScPD/50+Jm/Rn7leB2uIHHKE83N4oKvAnPL/3GG16ZBMexv3z
6bS4GcmWKlt/jahMZKtW4pX81Refzc3DHYclcjqZyTooaCQcgaxiAAcETUgVmJwN
I7O0g6Dp/A5euPneGsYgWwevFn79sJMuxwSQGbxXUW5+6MWLf23GEQ6IGREiBlrL
TCn6ppWbX+9eKTuwiPTEyJi88n9TQDj7xlH+VPCyzmbdoOPelDIKhey7/c56IbHH
qrSHCKmmGDz8YjctNXrvUWxWy1CgBbLjodT4CYZPWBhOq32hQfV0xWgYAnl9z6FA
PEIKQAFgEunDAeMnexTY7W6agXiy0LAvKZgcU0x4L96qwjExtnBlKD7kWooG9ZdW
nmrFUUOcRkwuhiWKE+ohRzD5/gtZhL0/dssiMBfnsQEWPttE6v8G4/Z2ifU0uw+w
VtWr/XYd5ClpoYlB9sW22OodJjhhsn99iX5TFsTLQvdAHAUgPPNb6UtQ+kR0yEXE
O8a08xCuLQRBD8UTiYJIktwOfBW8JESZhZjWkCdVAt9TMWkVvmbdftpV68x9izWM
nZNM3Xj7fLrFbTafdeks3WNa8YKkWqSyxcOX82Z7DA/w4XjQfUytrjnIZJ9/WANE
1smJRRzpBYCKIXOCpYovmLTXjg9vJ8SLiPFgZIpf6IpOKBA+ITAnISRqdSKHkqh1
FnhaaqNlqIEtgiW75A4OWyBfQbE/jjPP8HcWGQMf80PXgT+e4GcH/JOB/1RKFNet
39ytaqtZ6Wl3nlPYOQt/IJFQW2yIzJyyk1n5mGI7jmvC56DZFemgx6IJrYDaxWeN
J6mOWNVhny000M2eiVMj3oMECfl1Ojk3dUhRW3+5cs1lfqGwq7XtD8q7coOGjaA1
j64cpSXFdGu/EXZ6ooZpNpP7izSaR/cFhPIFdqbrUIma0j0Ibr2w5+xGT5j6bSrR
hHCJG6L2+FK/n1J/FulcqekMvsyXYyKY3sejayo/Pp4=
`protect END_PROTECTED
