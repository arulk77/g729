`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu477N8R5bHIBYvjSa5kU6vbY+1Zh8WDoQOpGTuVNVXmEa
j3gAp3GBsZqz1+UUdMANzJmMyzeIsFvB3kXJLEMw9oTbI/A/JOpiGoZbqlImHmk2
hZwc8bTcaOdR9oMCJruDKmQmhaQxaLxTaYEhDT0sQnZb1CrsG173zVtOrrFqwoOl
7DMLwoQuWnuMeymE/mrFPRA9pO3kpCdM1GEGnbPFPGs=
`protect END_PROTECTED
