`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8h8s1PGh2G1t29TaFLaevcSN+D3yd+QKx2FjZa/Ez7Z
qM+fcTbekSLKbnh4J9ZM5CwzhuGYg9tiyik5vqbg+AxLbwNZmU2E2CFUNpAtpElt
0qEmzQYxr6MTpfOwD9octrEhzlEzkZPlkRh1WL6Z+LgfMKYJtGPr4JniY1LOpX+K
Z4JTrG0sZ0YyTV+8nX0S52IfbWDMRNRa+1lSbYAgefhwnBh1v5gH+HKZ66nRan3v
HxFWQYCghoPQM7RQWRUNAahlIfwxdvLgMVYmB5+FSIOccwxCs2xgkXULZ2+U+qyE
jZ0FnBDVxA8fEFMsKmZswV9UdTM1avZ/AZ6Iy0vQYA7X+6qpumAx25OYQJYzJ/QA
5LH9oBUvbfRSrq/tjWxzzxZuQlbPOC5/JruUoQeYsRuRD4cvSxYGsf7wC5tyFZKn
J91OerZp5fTmmwOVi3uTzv3cY59TWKLxndZlDy8PJr15vzxEM+TngMqz830jLKDC
YaAiVnYlQTfr6wJt6u0QNB6mQw13ZR6rmMN4guFXfjPiUfgi9fqbi+lsFFw8aopw
YZvx7jB9Rmk4BWGWtddMg63WecNI34aZspxXQH5wYwnpiMTs8mKvRdWmHgY0T4/v
O+SrCsLFPc5XqJNQ+ZvVuT1Pp4TmzrQYvo7HqAjTMK+++w9ph4hQncSgKn6DUmrP
K/2VAh389b9PnnPUCQXBdXY9Rp1ib7DvROGBQNMzHlCGLah5zVxaXeo7WUcyjcju
V3hjlEAHkHVAem1K/WEDZaK31Lcubk+pev3EWqV2VCSL0n6tTdL4UcZni1tnF5Q2
qVkeQW7bQlmUqmIQXEs4rA==
`protect END_PROTECTED
