`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNtFu4gCl/bstm4B4zKcwsNkc00TnBt4qaY97Ir1oKBo
oM45YfBKxdM0ZrlBKrg2Fnr8iBu0TWboZZOQP9lX6GFPaqq+m8YBxbfTZy99mYJI
XSsQBg1eq7MlT1I8wp7blimjLAAqbd6+WyiBjltd69dcTtaP/Epz2bG7YH4F+r+F
4WIiIpsKrpNppvQ7U+i6MQ==
`protect END_PROTECTED
