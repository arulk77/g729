`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GON+rsTuGG/WttqOqfTOh28qqzlu9L712vEvCWJ0JeFhtqCuU2jvDAagrDTQxkOJ
b7bXSIL4BOP3xgzXdR8v0JGKVZJa7EuBbSaWM57LCMQX82oXQZBbOBj7ByCstB40
dPPPbiKikaAr+ju/2GVl9cs5MTLGRgZaHtauAX2xpcvOTDSyFKDR57dyTyOFCpgD
Pqd/rDnv3z4UkOEjEd1XthG/B16Hkl60DnVUi28oS9koywn/FWjk1StGGRge9IEN
V7C2WYqkQ8KtBG9YH2uw403uAGcknT5Xnuo7J4Et0qM0Qk1TdFnzHAhOje5P12te
xbgjT/SYG11yJOf7eio1VcwLBabeyWYuDH6H7inkiW9uXPewv1EyY6EX3+eXNIEv
I09P9I5HX7NyWgcjxFFsaZYmSNte9D1hdQEIerRpM0YM0aAaC3Oe5LU8bM+9tvGA
0Oc9o8BBzVEjDkINjpDJxoWkFXDGEs2KvzyaJ05gSVdaUa7UJSAChSxfLZXT+sXh
GYktH7A/yRv4fJtB7LT4hKz1saaOuC+cByXOnlgNIrKTY+AsaUENFsj44D0swZjX
2xZT4AhPRXDJlBE9O+YYjcZuytqZJ99mozFTSx0SKYwbCZuR4KM9eQtbGwKZOe7Z
zn6u6BTDVtgLZIi1EdGGuYbRk+RWY0gvAe9JUtnH8MMDPPCwl/gXYcSmxIq4vTAS
qPyX1C0kXT7cT6RrpDAxQSuzHr4DncMzF31VuuIn6rRw4Dr/ZIJJhRiE2XFvTrH7
HTeOdJbJ5Zje92DeErZLFbRBMS+ofNz7/IpVAnGjxnE4N8q55ajKaM+bmjQ/2QsF
VWwNw8Iu2aCW+QTDe7cTx88u4Y4FOTAA+INDDVBIdXCzmgeGm8RhD+4eSc7L+Equ
BHE/cW+CnfHldjIYkWa7FtRYyAA2uttTvYLyJXdVIEr80sbejNz+sONPhcygor4/
AVOE/sIj9kn8xa5UdeZ5i3inLWDUaNfp+2fRls8aAeJW0IMKDYAlFNIeoF4wPhMD
ZYd5JvPc8iQZDo9lp1aioA4X6pCC9lSfLmoXRfSrSrHKJjDhLpyenVyhvO30xcvC
TyWqVAUQ5+LCSJtC2vffHjoQ6fAklrH3hK2cI3yiiXZO6NZSNwA+kOCPvY1JOp/d
LRmdbnVjRGMttPVAglPjkAvO81zNyDj5a6Deyf7kcQJ4CBGRg1XPYGCQkpnQCaas
zd7LXT/ie4oiif2fwHK6QZEO78+iig+G4cY+2SA7Xz/cE6tb85hPa5pxxmzOLFqP
JxqX0fjNNFrPB9/SoXSaUSSZ+SGjIKr4fsZoFn0KVEp+3hUivlOY/mRXsBgKuEux
ban1nTRtqH0Ip7H+k6NujbL3t4FEx8HcgSm8fkmjhQ4hF59yig1LtYUppbBxLfVJ
cwW9i8i83ubX4lRz0FdNYsOMQE0o8q2mGxQY3PrixI3iFDVTVzPyXF2c26mcnPmT
5I4WZoEqsept1sRnc5lk8hautVbk14NymdvVrCerKshRe/Jt/KvCwoJQPvUBxK7L
+rEla5ipQ9N4sFVc+PYsJUvMfkBEFv2lwPZJAPTYjH3bKsndfIqiiw0pyQL7f40S
TgGX5GQ/Ln9zeQrdARLzqNITzfxop0SxOeC8cu5K5jgdj8qnTOhnTpK9toIYT52Z
s+HuZqHeW+1q3BG+yqQwdtP//Q39z112HgwYEBTklliZmgkwe9gPQHmnUfi9QJrR
hbIbzogfUNMzDhh9kx9E0waFpMxe7n4BaryVVUBQwMQgSDjiqA8UtE2zQiGbT1Cq
zZ/4DTfXc7whuB9MGKCMlHsMu7sQD1ZS8gm+9YjPzqemHyXbd814z1LjBqZDlkQW
hRzvub1VRkiH50DwC7zINAOoGjDDOWd/o51UdYcEIVJhLqiEIKr+D1mcRnaeXeoN
Q0f0oUkeWnYXI14XT7FPi2cgPhOyABgV/RJiy5QD8UZc0ta59qjsZVyiOV4pDN1G
1mG8dYLqHaQJQzVgMsLQDCP2bMsmaPEXxrXKDHcz6FB9vZDFQnhQikodrggpj/+X
wgVKhxGncVpG8Vm34jx2PPIhIIaACNvuNco4DCduvLd9hWZEvy8hhY/FMx5+PWtq
KY+MtbFeybZEAUlOh+9ftZgwemk62kjOuM8cimqlH/sCakWvGjdH2J8aCRvBCvjl
kq2CJY6tnO+QOK4tTywNTCZq+PXZIOcncAwztHRY83YY+VCrPbFU5Hv8PfX1zfgo
Qn19L8zgZt61vtWmubi1J3Zsh5P0R84NiO2IFvuH9UODbEIlzsMWtrLQsGSsj3ca
Z6Skf7Q4GJQaPSZl4RV2zA==
`protect END_PROTECTED
