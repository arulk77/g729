`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Cxkrq/4wTfFDlY8uYopYwZPonmKCtKBwpHoKPeL3L/gHsjgxZdTRyUux6WIBfrao
90GD1CgBTwpOc4sWjtUNA2mWd/YaAAH+oTxFaYKHgVwqw4v+UEH7Ol8n+zvmckKr
TGWXq8pcWg9eJpQoQME1AZFlbROHHX8UXe2cqXdSK16y9JVje0ut4VA0ySivtZUf
Jwgoa74bZVjnpbCSRXtutyFu83Iao0qELITJRumFc/G36Ylu/WTeq3dnoKytyl05
OvZZ8IIZ9DJBLVX9l8gSNUTipLLpKITCL+wRyQXORihtEbqp2d8nsMGgNlvTmmAm
+GWC9Ufv0LCjtf2gaiPuRL1IElVYEhOe/eCDzn0oPvWH0wKxjZtuCHaepwz/1Bey
CtHR9hepC9ohcBK2NPOf7Y7wZik/9i647Y6wYY2hEUHikXXn8PBVdv1RnIMUQNby
OP3SNiLzLlOQlkZl9/6aqGCHh8qhhXho4VTMgUJ9jKLV2uDHNMYmtGaXK9efV5P3
s9nyfCbst1T9pjvB+UAI/YPcOlSBAaYdz9+Uvu1qPbXm8bvlqwh2JeNrvpNc/jr+
Nfv5GmbT7nfbFFD67V3ku67bQXpis+E8BRb8WZ3fyhD34v68KO9ZTm2GP+Rcv91B
qpZkXI2ITr+9cEKQwY1q1pk5mzkE4VpNFQdR+/hYGqigNlWwPyFIZYgbJu6fFGsQ
fsZ2+l+RrE8/ygXxmgwb+Iyw4GDqAJR0nxjKYgCnnNlh1fCG4XXBUNT9S5kL3PVW
`protect END_PROTECTED
