`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIUCb1ekjY6VJtvQldEXUsZoHb4B3YRBa/RhHNQ1+Rwd
9MyS5jRIGVSpF3CTT50UYNusa4+KmzpkHy60KYHgAanBvf8oXswTvbwo2B/S1N4Q
I1rEbdQZIMbXRDATpc9L2+dIFTQhbhSm/8ryPWM/7eUkTUPY8Ys5uzRlVtrULeaK
oIC7ze3MmHw7yZGNTNqL0z2VL2cRlENIX01A6IJ+FvUAykMyQph3m9tUeWett/aC
RMbF3Dn3xn4CGx+HDWzzgwf7LKA1Y/212ZugIQ28qfrip/MgPmyrqdcxrWS5/Gcu
7Em3HWEXdRExbeSbvs01hQ==
`protect END_PROTECTED
