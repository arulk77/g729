`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aYSQHTXPA3PPq6L03Vpr7GcB8QenubTwseVAa1mTaLid
A0NZkOhC8vrEX58oFpisT83MPfTcD3WlyGOOGd7i6BBzUAxykLG979+NeV+y6R4B
tmWMoyaeXaSqTeBt+9s8zduIQgYeACoklk1kQP+qhN96FE/6Oli+ocFTKdzOJ4Zg
GPuRc/A3judFNHT/wbjz0ecuLQny9Sz/2e4R7zMD4zm/BAoHZtSbEivfmSv3EtUJ
6mBdoxk0Hyrhm+XXpfAHKKUJQkllnRe/std8A4X253AI5mYDtjY0Oo08ybLC65YA
hG4pgyPzxOAqBpY0V9VXpCPuFaNmNMeuGb8kNd2QDbz+SszfA3xh/I9rYIMWLGhJ
UbEE5VFgU5EBP0Lg4SVlyC0Neg8/Pu5QC1vw27wnqudVmxG9rnBctMaD3dmLHrYF
Ar4IxC7YRmsTwr3OUCANKyN9S3vSyu/xr3/YsZ+H4VS/aLoAz2ByRR+LAWG3FG1Z
tiTOnqzQUTMQVg1/GizAB3VW0zg40Oonny8xzJ+IUkec6U9n0TTatgbInfbMm9sJ
oTU3sQ0n+BPu1WqSxsMvxZsEttvHFQ/Mh9O9CtJZu9El+Bbt1fojVyUv0Qjr4rag
Oeic3cqJc0h3EMVteReSZ6OUMqN+8ZP6rg3BqAeK6kGRGrZR11BtTpUzYjnDGYz+
BYugApDJ4xuDSPIrlMmAHbLqK6owazcBNsFI9wQ2K/7+B3SQLmp5OAdnMUg5nXIO
nwb3TDiZ8tSmq4ozEdkfYFyEbSZOs6PC9W/VXdf+bCsjiSOFFPP39uMF4Kk5dycO
Ndn1SFUszd+dLUkkTdqt6atvtUMrTq7n/Xleq9PKUbzCRp1CWtlPKMULsp5Hw6/C
WJ7IpbuTJKd9UPyGElL+3+rKXE5I/rVeP9jS1TFmjvbUS+lU1IL+ony+BWidVB7P
YPaYcBWywSIOLEx8b9os75IKnqxzU75zPvEEwK++oz6rSRuWH3mckQ1sCeJBVlfM
Y/fSqtWdJANs5SpODdD5j/MmiBDGl64anVcepb84woB17koBBsd0hcnHPG97s7g/
PdN/uFzOLcJzYeBUjd3t5a5GBynCWUsQjy7yb2xHT4AN7wP6h3qQtI6pSuD5b8t9
Y45K3wENfnzGJq8w2Vrl8HdS2U9VsgAFH2+fdCWfzptPe/RT4nnJc7DfSnsxp13z
wJ+PKqJDYYO6WMJTqewPgg58q/QLF5AYC2VqAcIZ6g8lx4tV6DHcikIj/NK4qml4
oyn74LcMW5MM+W/VhhCQAz5EN7GT3E/aYRIEBLjUuf+8xXlDuK2LhelFiREnPn5q
8+P5yFH0NevKu6WeTTTH/+wZsNBr2d2wM72irpd4i6zkBXU+cXVB8GgSUx+G4QWQ
D5KfKL3YhQNAl0fGcO2kvWw0pvl5BOlr45r4o6rrGkF9GJtFBNXJFycGpDSFqefd
EuJp8i1vLfpESUUaiHf4wdT1lfqb+8A1VozjvqJ1yDgps2+yGrVQ9/wMhrtsKpdJ
WpuQbV6OO0pP4/EHtVmNdfJorDdgtUOynugnhJykX8Au+dmbX9VTB2DA7zspZFKU
JUHhForXj8Jj5N1VdLdBEHw4lfomViV7QFSb9DmEuYfvNdxQgmX+LFljU38qrWr1
D6bJYATNTsjFGFEqNPQL+snxCj9yJ6A8RyM3Pn9MAgRR9YBUBhup5pyv3kGPTj7D
dS1WUtqd10lmO9i4bw4oakdAZZ0EYoe4UFsMITu95Lhrd7Gb7aX7Res6PAYMj7ea
0m9nlXQnd1ZXckr3NsWvyyrwYtIOL0Eve3Zet4N0xLb2q0I0oANlrddObhUf1t+w
KWGXT6duUMUdIIqEkH39qX3hMr7f9v9RVovfElACZDiH3GTJ8ecFukPdQPihhlAO
rnZ72SJ1NvXjg8BQ8gNeKRKaMUPtJP3u+tq15y64CYHc0f2T5Ky9lkUdUL9KbimB
NGXVnG0vJhX1O2b7o1NvPTdzhPJpfDvZdU0zNKi+WgMyg0E8eGEwnP5GlRahN6BB
R8b5iWlrUWOQceWh3eiGESaQ1lAM+WcXcL8xLwPUYCJtozWbUvfSJ+UjUuZROZtN
GPlZ7f7wZ5IsWqOgaBfzVqpmfmerO1ZHseGGNAJ5AUdx3Df3bnvBnb2cSdXHq03B
gFauHwDC/+1OC1wRybW2w7uSyZzK3Q0J+7+t0sGyVRiq/Vk+vjlxs+BUNcnzh4r4
jnHszK9EeVM2iqBnyru2kC8n0TMietANojnvrE7LQ/00PWv63894EjKuxZ/ZNqnr
vExwRRgPDI/cG6vhB6ocWp0X+ZFRWnsi7NrJ+N5wIM2v2XbloL0g8m94I/1FNqHY
8G3gJHdIw+lhNHWyTiRsAgfL5UAopB9F6HSKCYvwi8nRO499cK0gqlK73qt/rYsm
DiVzS0vKy0Mg/XpMLWknlG+nC//eM/2wrYjrBPVVEm5vuxcUBRP34SNtzgslFnln
w+VFOhUAUDgS6mFAgC5KQuWEnHIWfV7OaCg8toilJ6ataWJLs4jL3SZJ2F5imDY+
u18zVdXMMeR7Lz8FIag7yew1XZwh9gIghLNZBqnyIvWLpEcaMHoLUyGkZ7atEVOp
UCtk5mgTTpQgw93/aEon5xz2XV7shuZDNB2dlTD/PzSwddXWWa1piX1bJ3mvGYZ5
NPXYNk8qqwjCfB12r5DOKsNMs5Fl0Odh1Y/RNEh9BD70Ohk8Q3fSsl+MER4TyNjt
IynWQjWufArGrXswGupi6+wCJ1nSvMGEU5Pf150F6UPNYyHuEF2DTpddQJCtboo6
+xtIYrDyS5cVZDSVSnrDE9ukiJEIkVe2tpHhwzlwann4DVZck3HS/8Maz5AmDMOi
eVWyfqZPeyVYa1Ug6EXTZdCxIwHgn4LUBEuudSjzj040HqISd+PcEaKXNiTIyaMB
jCcXsRuXePWEbMQfram15haSP2RIKxnmHW/K+3a5rVmuVfOErwlCzHLdskhs5siD
7t/5ySYUR6bPRAWaqUHkuN7kQMOVSHrlqjqNfohzeGNi7xb2WCt2Xpkp2zfL9788
FMRrlAdeTQW1uFmvtieSWs+y6AVbHHuyZ9BpKxFlgMF9wbanLRbqvbDRANzMzD+b
V771cCYAZdAktdnU3mDXj7BeHpZsjanOjA3dQdfwunzC/G5dxQObf5iRF0frm0z0
q773+V7UEeeDrZ7/q5ArTkqYs03y0ezjxToALH3NPFI6SfJEN3YHwW0AZfP24+n9
iTL3rhKmPwpHHG9NPy2B8SuWs481vSSmCA14vo7uN/HyCBOcA6qCb7lyj9sLgn1y
ONKrLtgOJeSQrUMG8Xw5+bUl3zhR322t87mi6y8VtCUi/qfaVRcARgSIrDBUOORi
SoXt6RSYB7GdAidW5N/zU1xD7INSTdI+z1E6Inye6DxAxBizs/xrWa0/sLoLbJBU
d5dTEzg+d4GBJ29pPlVdhe7aeCSoIwpBZlB2GnB3Ie8=
`protect END_PROTECTED
