`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHbZXuF2vX5lllPpvhSL88OPZCZXzyL+FmwDolSBgkOZ
e3TBktgjA2YSaO2HBqgHIlC19qmbEds3MLHlw84U6vq9q+lcw3mTsbultxjfAMOe
yP3Pj1gB07UUQjaMD+qS56VfQfKLvHiZczG3CQj9+Y7w3TgWgg5Uu/D1/Q17DDr0
sHZKjJ7J66itBhpjgNxA6mvJaW77ERlvHd46mMqwre8OeRRp05ke6BqXfXSDVU1y
aCfyIReLRoB/GHTwKAYBfeDkSE7+7Ndg+TGwVceM1CeuW/nTKiiuri1XnWPg8UUc
0CDgCo4okeztk3CnvmqiA40e1aI+UB4TtLBx7iQNse1A4wBC8RTDkOTQn3Q7EC3Q
dJCuab2Zu7QRNBi2O8uR6qdRtZNM/hAEdJ6nYykKzD/DiH7M9u/BptMPua4Sf9bD
Jyf1ixoL1pRC85k2AllcUic4No1dzhArb9kg/fzW9dHqmDPJNH6fqzoP5SQV64Hn
pgK3IUwbuApZagpHgPIo+USUCpiVT2einaD5AElnY8DYXqsIyCVMJPkBTIgazGxs
`protect END_PROTECTED
