`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMzwbSgUbl3oc9EOzeG6FwV0LUpJ9yUz7w2gZyY5Ng85
X0XPWDrmgqRI8e9oOHTOm1yYKyqB2P+AGlQxUgkpQPFjDPIZoL21HAn8DeXy0rH7
gWg7O1W8y2uVGtoWX9UGGZWOKBYSHNF4mfcr7ANYi/WpYLvZ3OfsrQe0oqYfacm1
l+D5oLgSDfeXXccCZfZ3gUgUMX7KYgtdzuQF+wCTNBW0yYh4tvvN2DWFVqR5be8w
hn99AQAmP8z5ihzkdMH/aEJsFUSQ0zvUF/CWGfBldujGvafChUd1Hmc43kHqCfMV
ULP9bz/Ok3kd79ZEpqb7Trsang6Ip3/tb5qasX30hnnOQmwLkmEb7HD9914PZxdG
CMHcL9MmZP7tSILZVJARCjBfzGHmEAmU7/cJf7x7rZrdbCVJqDrWSS3jPD0pMixG
6UCIaQq5sIV5erc4XMihpgDV25PBP7GBl8KubyB13VxvTqPSPdTJGFk76VLjD/QT
`protect END_PROTECTED
