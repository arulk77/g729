`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveINevAUPWmtEpNiA/OWrcbgzFZXCRtNar0RyZJYRL12W
CjBZbtpNdQegfEvgvxfV7NZcVoLaTTaBK6uoUh/vBOy6Pa9GFC0+Iv+QjdIg73eP
JGBUFw4z0NLSOWMEcH791Wxe5XsWRRX0ShHRQKTGImbhyYgPkRytQnL2YRGo/oRt
f8KKciA2dG1HE9FtX+90MoEAss6CxqK2dfq4AKrE1PgURp6nndMJ3ntCPDp6CfZ9
uQrZSNrkK5kvVyIjR542dToH/o+2CGl3KO9KSxI+j+PTV9E/gke2dnhNqJUmnY51
splLnZz4+8gNLRKRdVIm42FgMZ1vaVp6JJgXF+irvjvYEBXaLTe75puRGnogGGn4
wRj4+5BP8YIauWZH49cIF5RnIIBEU9qDkPKyohAlenUE8CQI9RZo32/u7JjCTy5S
nkHq6WtJYbdAvonTqKrgunOMVkqBNfATrQ+yXkpqi3JbRTHmvy7XytGOeDu4HsmT
tlyohmpmnAM5yXiR+FYb8mPUsfmg2YbRJrjikBK4lEQnmakxzBhGCj6ZeZ7gJQ4O
4EyeL6jF5xLwNyD2SUbeFdodgKLpJguZvCQqvEhS2JeFDstzuzwd3KAyn4uHpzr9
`protect END_PROTECTED
