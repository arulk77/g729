`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43hJ/JkOAnHEKt4Ozydu7aLfjQ5sufv8dD2tardlqNRV
87zzwLmG1OriHlvd6nW5eHXc0m7UcjoW+HNJ5PgN8rfLWQB/LuYQvR9ul9ClElvi
XhMjPhe78yfMU/HNbpUB6gu70MRxx/kH/BAXlpj7I4pJQg5uPvL5K7CfRyYDJOH7
Ac7vgwMjdCa0r0LjJ7/XzMK4whrQciAsfsPtdwMlJhY8s+WeR+Zzy0TNpjh4skSw
JjG95xCpAH2XVfsFBWyU0ytHEsct73ZyGUVgVRfW0M3xomEtUe6E7j3EaVcsi+lI
fSggWyRy8CduWsN5Da+dSvx7APScCV8zml3T1tizJuVNQM8td+e99DgwPOKD1/kT
+RC42css5Pe26WOQWfRmZfqP8uf195RxzEeXHjHU3JfpYRuL71HymsfnmTTU+5qK
wGo/fJCgkbxSr/bNYvHYLKyH0nabwzAIIOuc5SLIm5Q8sIsUGNWXxkl8JcTXe3KY
`protect END_PROTECTED
