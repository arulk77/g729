`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMRr1a7XmuEQF4fVH8rUU+ua7C0eCnYlBwZs6tcXBLyo
m257/LFL7U+RK42QarmsUXp8wSaDFDzHpxQPKRft98Nj/xGyvxjgonMvGHEQuijo
LNm4yDq3Q0mT4v8TOaWIBlz0P95S8ZRdHHdWtkm6UGF3Us4t3vAm0rKaUMTlkgl7
pMLyCsT2jeDZs8Z56NUWUpoDJLfJzydNQHXjFKOZtDveWT44BaUAmZk8QSfPuOU7
LI4VJJ5btuHwG0sdv2k3KQ==
`protect END_PROTECTED
