`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43kKKprGjsP3cE06sXFGXgvaBpmoDY4bB/qfdoivhKVJ
HQJMSu+QjlErEDbTiDjmOSIRpW8wyGB3WdARu7bT1zRw3rcJfPlkSTIIkrx2BX1m
2Cy2DjyLpq2Ci4bJZJ++ZLg7D8smt96/E3BaY/RvHuww8be5Dpgnha781vvC84wF
bIb+65s8XYq3s9mjrxZvS6njkPNWhKG3mBzrk5rhry+PmwBhqqteOh/YB/87TZyz
1rrLCFDy9G4Y2E/iIn/z8GsIhrkHEgEd3LMxDfvWdRW5x9flvu8lmsBJmtRWOWjX
ibccCQyLffWLT5Jo3JW9HA==
`protect END_PROTECTED
