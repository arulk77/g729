`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAVP/vTG+l4xklO27CUx2Ti5rz+xCpArqxib+gaUl94X
59QI/q7ODQq75Igll3Npborsizi4M/8+AvI0teJ100qn9mKeNn1G0PRMKfhKdfiU
ejZmgG9UxUi/EzB8oNi9X+iFzc+yaarvQnqXDd4cguK2KZgimWQNMr+ECM3rD0y+
lcXtb06xTelwT2yl8Eym5MFDY67dHSGA1jbI+/M6QkhYK6yZLbE0O8ix7p1vx8AP
`protect END_PROTECTED
