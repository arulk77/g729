`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGP4Ma7PPQU2/t4Jzrw/md9v0CKrSsbihe2Bi6BrRzU0
eEKriYRhGie40VKcCWlO5ujKVf3X2pzQ4KFYMBDqKC90VFzDLntYTnGwaZ/o+w/K
mE2FgGh534/NnvQeVgIIS+3cFeD3dzBKpKNGK2sMTe91EkPU21QVEGpTzrUYHw9c
yQY95WItoH9z26Cj9kD+2l14ZgW22p68P32IYSovvbkCG8QK6UDXEHvZjSNWQoKc
`protect END_PROTECTED
