`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveALxWoHTMK9KX+gxokc9GcannrWDt6gs9yoWl5514V0j
psFD4DcOfqbVEJEYSvqkr2SNAzv1uGToWyoCJBRtZBsijKssQnzFaJQ44GQFnq1B
OIguQhcHn0TRrBDMYSDS8uHDPMDe2DV7BBHRoeu9oiMPwBwO4vSQI+0UEVa2q/hX
RtWC3KfuONI26Q34/JNMWSgGTm9dOgpQ8x+W1j0E6ROcmSVUDpK3OWO5ruIhTO77
9Cz1dwkUk09Rzq8bisy+tfT9FI8xt1sTO9Im0hHQ07q4oZjlncx8r4Eu4IGp5p00
QsFobl74acYW8sPGe1phppx6Ol8IBt6jMXp8nMcFSDNxaRaa5EF+d1E+Ox2VIKPF
dAOrh4rvp31sYm0WDqXoLUW5lkxdDazLZlE8JyOKEHjMEMc/AbbgEcfkJSmXHw+w
`protect END_PROTECTED
