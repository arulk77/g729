`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4y5PEQC3iMionc2VHE0Vt0abM0UO1RkTQChSXFxdIZUA
HvuHkKnK5dn+oBig4bVkUmlS/ChW4jpGBPHhuJ7hK6Sl6YVW5KqHnBOFjP9FbB8N
KurzBOdUL9Q5tkTNtg1Y/wsgJJTFoX3u2H6LeLfykFNiIo2YrcR+sDtS/S3iSFz6
TSF11op4Esgj03GIHyf7BkEcl7Aer/Wg6+Mly9NKUf3i8qVnEXrAyRr/tYkTy7jo
KLzoQcYmkiJFP+yAVy/y3AuvGmy2iHn/s/uZ72DU4LXbgWAHpIv18dsNVQvqcSWX
dL5024yUWCqkjQ/Lhuip9w==
`protect END_PROTECTED
