`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNDTCQtOvduw9CNAuNsaA/fKOjwoNQsBGhTI1XK4DyqD
ULq1wbaBoCT/wvh3Fkd3sRsDnH+izYI+8Bk/5RULsU8wCedTxTd99mtPOMNW7HCM
9qnTsTbnx7u/0WhLzSXFmoW4IG1CmaHsMxtKAkB/jBBIN5gCqJfGczYfRiIYNUBE
B6Vl7ZdzTfNdZCekj1hgGh5D+oK7rJ8hOZ8xKk27++ivmiOc8BwVi6Id/3GdmHQb
`protect END_PROTECTED
