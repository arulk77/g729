`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43qk0iUpEr0Fc1jJsBNPMXq6Yl5Bg+TsPbyf0grb/wdm
EQyR66ijoK+11LOQTEa1qkW8/BUVvxKBn/iqyfkMOhkWZQArlrO3ejVUB5yqEyqq
+dzpgcSboeP/6vm7B9+faG1LUjYhR6qVpHpzzjDelpVHYwq+CVV5v43Snljgt4GW
ckHBd0c8lxC8DxedSe0HQw5hQy4apArNw2IDeyTe2BEnTUMPujyszERwZwOEWTr6
tBMVgtGpviac04OU8+4GDiBiBap9CayjsYdVTkIeR2w=
`protect END_PROTECTED
