`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOe+13lMy/vbPsuIDtt/PyqtdrV1xYiXfJC18KzvV5Gg
fqR+FWN6y6K3iC7WXRi7SbqXgAgkwTp9JDpEpLUb0x7aICX27ZfECnUmg513JbzP
ZX3krrn6rQikhYWIEOq4H5aCjb3Seym3nRcThXzArTlEyoijenWGDo27LRpd3TeX
smglwvki5A489N4lGox8ZtzQp2ol6zjR37fgFl/9cJU22OHmijcIUDyrXsi94dv6
V88b9A5fO5EfGAACPzwuSJaMdQonMIXVBlXC+dHXu8MN6u9kNRZC0XAeZkRkKMuO
IaftBu5a9v8yKna31qi6/w==
`protect END_PROTECTED
