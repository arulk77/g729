`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePbQuoCrqmyRbDlCm/Gcrm9NrpOveKF6kyCKoS/Xu+qP
RRHIV2BH0uEXv48LMU7CqZLDA+dq3fkElUd3EiFwwK9nVDkfowGyQmVcPzO73yzb
epOaYFFeXmYS/7Ta4zlSBQJ9BDZsW7PdQ/n9mEicyQfbPtZ2N2TuAnJYnT/S7Ni9
qXG3yhk7XI/VEQRc/6wJ/e4ZgZGN2l2uI72KbuiZY2SkF1HmfIxVMxqH6KLAyvI3
JLGnUoKbc6oVkg9aLLvKCc+94lrEG7Y90XriVdwH9AkerFOxeDA3KHCyehmb3sAc
eyDunNfw4ZTWMW/EHg5UtOojI4c+swZLmIh0kxTCWnUIzfqovzyUzTGtjHOw0Y1A
dTIVQCbL3h7okF7vQfKR03U8aBjK19PPwFB9ccHfEc7k9Wzk7IqR/b4UMeFCd6Io
49O70XfapFOSdj8fBpghSP6Y++iIvYEFUUG3k0lxxsFMlYlNhukdngTUU4+U3JLT
7Sb2KRcZ/BNqYljhazmkBlIK6hY90FWTUq0Zf/sA4cnbY0JVsVxsB+r4SOCdPHkC
`protect END_PROTECTED
