`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xmqX1Wlh0OuOTSZ9hCG+UEHLfQjVQQXLyX0wd6mD9HM
zzZch6Ri8aA4Hx16LhSW7Cvw5tX86bH7BLv+hsBElz/l8+NtFH6eKl4gb9R4DHyr
tR66n3CjnM625NQVZoTyYY1kvmyJUMjSfI4QUCsmpYnNOCaGa5sYQqFTDAUC2j2n
uLiFaWRRsKuIYbBopuIl4ZdFSeVGS5Iqd2VXI/IRvhQ=
`protect END_PROTECTED
