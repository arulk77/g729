`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAQSXfGNB42Np81l4W6tQjnfwn5obBZ1+ujXabte0rpS7
0YsY72YKDCGiRaqbD3YroJq2CbnfuVqAEBQv/q5s0iAYHRpklC4HTrsl8ZJNkk+e
tzM8llX6fl+H2RRFbnk5vMat+kvQDPAjMDwlYC0uq6tEhoi6UHIRns8cxjWyL4sg
1LOBP+fKU1qFj6kJQpkVwFFQxiTVMLmqqtfpOF7YvRyNXv5lSQ4wiCrL2+lN36sW
pYm7/BDa9StMFr6PY6Puylxia2qns1RGEXiFjGzSyaBcSSvbdHFw7Gy6pPiUsqFC
M52vf4VfCSYXY50KNO4THYMHvNVU52hUASXfx1IVSOrWCDGpy30MIyIOkG4sMle3
lmSKofPBUcYzoZG9BXMYJABCJWttMisMEvnrlePaGkBz17xmij0Tf1wrKoSAS8vt
+ehoismopV5D86ltlT/hqohHBjwtWHBlWeOdSydNDYvpaCPluyuZVz8ED8HJkuDl
XlGg8ulVfy4vAbMJgyhQ1GDcQjAPOd0g7OAlzYrTDdizRjR1XANjebMX9wvqFCkH
/5awzTfQDpj4V95a9rhl8G99aohZO5ybDlL2lDa0YX2FaUeuSZJxGuB2xv05fUOm
RdR/oyIwDj0A+YxQqEgvPh/ThtBeWKfc0Ac6LMYLWMsiMYLyezQyQsaALfkBXYt9
xmy5g+cOxRpWmSw5REaxlMgmmeq/mw8BJl1T32TMWOsX94ZVz7D8R3xzwy5p6aoW
hKNbjiW4fh/0W8Qx7xF0STnLuNKtL7znzUg89grs1owX5h+1kMm/+kYcxbZTb+PK
c+kgpt7GG5IlyPSn35sPjxZ3k8jAm8WO7nX4ex4hLMvyvwLqmd/TbrEJcU+v3Oyb
JwEJP7QTpejJ0Dzps2F+DPcqrZlekQpFT/+XpW5idRNRMM3qdWdM55QIL3nowIZC
2BKN3S1kOGU+P3qHQ6/pgMGazam7HovkYDo6SZ+k87yYqGcnXvv+E2kWtryHPh60
Rvenas9Db2CQxHFzMEyGVIqJrj9quUvCtFo7VkX6inSBvFN6iAuBCnx7MPFkhnZ+
oD2jQt9UeEO5M1+nBHDhrEkb0mPvFmRWMbV5A3nHxjEg/h7YKiIxaZy6ucRbjcCq
vTFrnGkRZ5okbusBJxN8If9rAP6M1CXK6Njs66K3ChSy1qoYWCR0Mb3TBIIUmn8/
vTdcMKnj4h6eEwyRbA3Q9jqAnycCIjlZ92+KQ90LjZIDcngU+EPq4+yXEZJgjBIM
GzZNGmGcKfVsNS90MCZN/i9iNFZItlmrVdtqbVEDt1jeiC0/RzNaZ3Np12FS8eE0
3J19XnD4QCWv5mBFY5T5sbY8YS4bGYsoMvp+Caa/i0xu9hJ298mwYHKDpOBpz/IO
fsxt+tbLfzT84RWwHh1i278erdfmClAOlWQ0RfL5z381HI5CkoUALhX8KFJ3NXh0
VLvmsYshz0SjaUzNYdRlXh+x08ealflqCqUyRa3TVGWGGDWI+sTXqEhxmN6I9GqM
ekpHUS6ayey5Zk1B8b4bujwPQXQuf3P1B/TWnGtekA+VVu7vlQ0kePcaAbyPq4eS
JO9uHMkGd7wSxSH6rRBOHfckwdHfE/5yMM4d3s8CPCTYtLhi2pkc6SC/wFPdbMa7
m2CRFWrg2Yy4VNVYdBk4OYFBBNrZctGMc9U7pKSrIonaZIU+7FphOjFPSJi+gfbQ
m55HmMgoRxCIIjAt4fR4ElFP42vMsZNvI+X0X1pwTk8nQ4dA/fNHhrP0jRxrhPRw
4AegxixQbpoAAff/v+Nyyua9TJ46wm1M0gLJswUyhADEHeJBLtv9QOof9OBlzglG
7LFWh4gwSs5r1rgay2JjQwxm1GqRTpxcpiRo3vMKURrEi+mxQI55FSk0UNB0sQNf
6t7bCSXJpR1yuQwBUsLVHitl1799q7UQOam95IqCDXZb+K3+DROHytIgR704CO0g
yBswE4OeOY5NgwnBxWhT80H9ZEVZTDuFpraWS5xe7CtdyG863UkStcHBoCuTxoCj
5RLVqXOcFyrip4JcGwt27ydG/INbE3nHB5naLFtR6vR67KKGMD0r51IK3rN9QwB0
IPhsluvUsZXa6g0Vao/AJb6EY6dji33psrMkLF8XglD57VaC/5ROohuojke+pN2c
VIIOiwTDqwpAKcPSTA7DMoMVdR2uF1Z6VILRXqXi59BdqnhT5zQc28x9oDDgvqC1
CgqqxWQWObKIDOMtGlswGrY2Qj75gEGq6sldJ9igPa02vsHJ4ZrPD4Bk52YZ0zc8
LHDgj1Kva1GqFYCSxSiI15SoSYbdmRQNnbifrExQVII8bwaHLx3000NvyaIOMf+t
WSYN+IHqTeEpCyuK5F3L78YfzO19w1qYIhR610ACHqA7rIck9EQsDh1F30IpCh+V
WO0HHcoRFEiqVy62/fYe3GvyvQVnDIca3bUT4TFaaMsofWBHSpZJmRyo4kwW78pw
ev7HprjN9VPHDm1z6TXEhwunAeH4fTxk20Jt16bAT9qYk8pYu1Keyl6r45peFACD
o4LI7WZoV9NzP4FiOdpVqcnyGNlxBLLqIQkTZd0ec1XEYBVZh0+aRfyEQWN2YzoH
mj0IwC6nyZtfa6++Tc22E4lqKxUrkSnlJxrdhDbsIOf6KZvjt7BdX5md+rHaNLfx
9zOoPqXNoN1omsbhYlUU0Dt1l80IhDtbL0NZ5cUocwlh8skVGcqJ2jSdQc9ADgUR
ze3BllCSvLkAVZH6vHhJLjTeNVA2eaaeOQCTw4mTr6JVj7OzSinTzY8iKF1KcSyh
W28Ws1EWXP9iPjZLYrIkaeRTwNuYzUDHExHke560ZJlcV4d++At4Np7tmu4iVv+L
tI1++WUF/pX+JjXOA+QoWkBk0hwgo/hADRjTTuOZANbNEjgdSAJL0hbjgSwQMS5+
hyQGeZ4jC0e4Wbes10DHe7LCVj6/LErsviX2K5JBAauCeJoiT1p48sEvi+hWoGMB
GGd4GeEURtGLT17wQoIJOvctWPY3OJeJ7fF4wK367uJlFbCaxw7FS3VOCzKKfjyO
sYT2/aFSeMFlWsJF9+FQGzjJy8lQpNxZyiEfstsKGE+XT4Jx8a6ydM0grozh/QAH
ynNmEQSe3Rpb+VO78QH/BqaUR9yC4lX4SdFz08qbeGDnp89qrMkIJ4XmvCIb/HJM
G6/2n05PBSMCkxwgubP1AgRIJB62UkELwxbfQr3j0WZ/iO/JTPGMoEPFuKsGSjHH
rrb4WCmrmgsRl0p5uFNP258il8zi1ioCbElcrKW5MofZrteZmH6wNiroeNwOj8Eq
iO+tvZ/G0saLuvWwDmUruTcbpq6QzakNj2neURi0tOg/hWsPHSgIRPhoans/xIa6
cpLhg7DXKsqPPff3+G5yckJxyhZRmbn9+RsEVXdPtMaE0qy9a356yU1MX8nxXQu6
4CrRzjuBKg9RL8DxE6e1ywqQaNB9wQjIUMl1Bqvc7rIt8AFgyMYVNjDZgrU/Fa5Z
J54IfkTUpdr3gVacSRVd0U0eOnikf2971uY8jQFnv3gHXbkGR0nGL0Dd5wzB6wij
hNx/onoPCDizyN3MtYf78AiemPd7rgx5agXv9g85AWI17ZZOJipDhx/9WiKPuLgR
9LkobenY/5tI50ncErgXHS4Ft5UCoArS5rWkLwaht3+PSPcCc6y7TXeAT4PQ2mCI
1wye2oyrfaFkcJmpMpyCUyO/qhdJXBwvone0q/RiWmcpLIS3mPmXUgRJEhHH2/Ik
jXg/B33KxjnJvEGjo2jO+0xYRj7aoYBwsmhERbdxHrOcvM/qhbttPylgXBCVJBbl
Q9cXe6qKP10xa7aVMy2XP1/jT1gyJNc/7GbOsCaT4C1nvf2NjXqFOU5LigajKkBB
u0RzugO9CK14/HYft+QlN/adlW/6ejvEoJDwRBippT4nygrA7XmUaDq1SWJcUJZ4
TYsJpEZxI1NbEBsdCwI4AFCNT3wb790asQaHMe9vffYMirlzSqt52zzem1XJt/FC
`protect END_PROTECTED
