`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
C9sI54IyUfxG/jrSW4zo4XpWnTCnzC2b4FpB91zClo0aHZFuPDZigjFmjcBdya5F
L0iwxnMYztGh4rCzxWumMjYUmfMEN0vFslDZqMJlj4c196Hs8WYBMgge4z0fv0Eo
B3/YiKPUZfdmyMecgO4LKdn6/01ccVzkpwmzeERDwYpEWKRX3WmRbCsW6IYq3CTz
1N6O9371zjAS60huoUKnIoWw6cioicKv5hDxgnfo3bs7QZjBIVyCwfpCwcwIiK3h
f6eD38cRVtArk+EgvTIE58aCw+gPZjYctZnAfcROWyA0P9MmRtdg5vvKsxhvJ3Hl
`protect END_PROTECTED
