`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49t0mJLN4SXNv/L+LERceR8uNuBl8eMrtW3OKlW/RRz+
e5PP8NoH+riH6AKu9Jq5GLZNjXWrqYjQdyrC0d8fvIt11pZWgiW8WxOGdkWL8j6H
v+uBcpTyvXn7WlLK1IU7AAQJNJBoeCLBZgb7ydjmkT0TpEzIZpMsCqHQOA6tHNRz
d+X5qSX4l+HqEqiaPmbA629tGAfV1X54sPzEsIVwSns=
`protect END_PROTECTED
