`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAMhwHcokcDD7eJYwAAl2mCr2v6zel8ZAj3bTJUpuQ5C
NHdzijhhe9b/VMyviQY5kGBVwMK5u/tWapvuXVeBcIU9jWXGidfG/EnM5XKEjw4Y
va2eu0uw2u2xqqzuB3O5trPUZJ/feWtOTCH+iDQyZtu+oP64V6vnrxLuxoMufTQX
RqAQO/rfUcbEm+ttcnizo7p2B3t9ekK1zAGNJwIiSFFqpW70VVhfZZz+G9G0BSJk
dDttUsI97FOT/uJ4vos42S8oKWhThc6mnlGVP06Mb7S6mEDw/hfLsl9+VxFZOGui
Wn8SQhccMnByXufVBiPS7B73EYfH1YfpH8GH43JphbXGIci+eX3d5F9xbb50QQXr
a6jYe5KgRsYRbLdgP2fZGbFqq1/dYI60FcfgbgUED3U=
`protect END_PROTECTED
