`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SaGv0mSe0nrP2R9tIkj4XGToJm6ixH88B1hlYEGHzsQH
co24an2WGGe5IYsh5Dspn/wFBewSFnbJr4QgC8hPntneNs87GvLuojTUQ7PNAbHL
l3OT13k4+Tsob0okmINmABAnOC4KQJsC19XT1HMuZwsGclz1JmuvQGIcMNQgC8do
8XPl+lSnEJ7BM87P4JUGENs7Xp1FIw0jl3cdgfBpYfMJiVuyr2v17SDx8D92LQhJ
JvpXH0NE7W/Ocm5j3ZFDX98JFtTjQgd4Qm98tgy7DpvNjRt6Sf2meQCeDUGUMZxW
pWDvZOPKATSlmtuJ7f54Obxnt34AMV+IzD8Igcjz1Q8FWqre13WkmZ+roJiBaD4T
UJP68rXAR4XB3MNLCTlBQjBLpNKagcfbsVOzMTAk2Q4u9Zfb/XYvQr/pCmno5L0y
Mvf8vUhSF3BP06RoYZjXG/ddNTDDZMahZV4RIzk2i4bveDepYy2EM6EoEZmx8RrN
W4dh32txwHXOTPwdQqzDcTgcNCCDfKYQXALbj5dy2mf+2tiksJ/EGa6We4XaAfq3
xChpMDpUuGt6xA+FaTMCA2ugQH5xevteRo0pBjOFMvKAeKXIWLV8/leq3nFu1IEv
22econQrDf/nBrzivX7ZwhNolBmvFW74kaCa96qz+iPoz0khh1i+9vwqzJCE35IE
lL051xuzx7zpbDqm7wdPxH30MlbEx6xV+XUsRgWBo1g/3sOypMndbanvFs33cs8z
4I/nLBHHjAU/9IZud0qZEToHUxA4ityaXfbXN709OIyJnW3C89k0uDpt1PtGln5b
TVwhAMc8jFpTaTpyeJkbxna/+GKw/e0S8XanEdGU0ok4n39VNUMYypVawnUAewlf
BM141400M3X3zhOXekGgSbzBo3LmYFfx7JHxu7oiK6HDSCiWaCTHwxLHKuu8kzgX
zVek1g+wkG5ElhdLh3pQo3dsoygyMHe25KriDCtBSlo=
`protect END_PROTECTED
