`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C/PNKHIMQb38X0rYDXsUo+8/kalTnNFFQDOdqakTi0mb
yQYDopmGpXfVZED5wOkvXzUAxgQI/bo3WIGZJhxeTobVHSynkTV9HBrjJH525a6T
AZW3iTeeymq77vh6qSjY9W7hiFffSDt8k3YN9yyPUvMNdBkJOtnUYIHMHs2o/Rvz
6nrScx6WwE2ORf8LYKwsp8ZTCo3sn4CmwddGRNuu8FT6vFZ445qUbog+dK5Iyqlc
/iqICp/Lo7Cmxz7xkb8BGMK5cTzgRji9COypBUAMpDCjR5AOY0bJhEgSbgvdv8fh
fLL7ebz9/qjaGaPrV1tDr5LoyeUJd2ZwMqLWF7Ke2+o6tztvuqCKhS2cVYPWFZw5
WUBsFj+y+BDpElC56TqPDDYoiBqaWxkCcFY25YWSgt3QXB8iob2zeD5yVGVFm3Ox
aQepgji5nw7n7HLRSsEmhgm5SLs/OY+VVQzBGOLgR1hdRPgcOnRdsdFpn7kgCHg1
TmQ0mKmR6LEovmcFMbyGnSwzpUU0xwhaHSW1rZidEB8WnpX7VUc/y6egQyKXwnk2
KS1MpOS8ZC4Su+iIjmujMvND6WkhK6Ted33Bzr6B3+ymg2OO+I9R/060zjGXKtkO
ZbTssqRsIrYEGl8Jye4sSXG7UTQvInrYmzYSYOiUc7IPI3jiGJn5UDuLX+KP33/C
fhqCuHbJ8e8ooAuC7OAxTS45kw4eZhKYsCywEm8pkWUHH0Sby6eyaLw1oWPzEz94
4qVMaQPG52uqF6D1fmFBTubGTMcVoK9v/qSXnhgJaEqv4ih4mzlJO71YEyYM0Uw+
/HclSD8GJU6tNh4yyKnQ57uv/pmw4YBGYuOkitgYwfnAonguPQ255VVdA56PCw1b
JHscxC1RJ6jQwz4T6PCTWZBB14Luq1mD/cGGGtBAnpcA3g/gjgiQivMUs8qRo4/k
3uaN8y6RFJpkxi+WfBH+qfHImJrzcL7PuWi8kVYNJQuqiwkZYYfISX27VKQdCpVt
Qw2q+oG8aVY04h6lD0183ZXvUxD4ijo0T27+qwe0eKUb7cInatgTITBMQ9l8Pc0A
HoKgwK6Q7VXi/WhdpG6pfJRCuYI6weTp6r2wbJp9wSD7JXGSVlSzzFx+GyXEaT8N
GL36AOEDoYoLkD3yHmCzCzfJ4jJEH7gY3CYRyjrOgufTb+InCyp9wc99YoUMMUrR
HPycnc2uRW5nRuklSjYO4kIvjlDHf8iKIGqtxfC3nvb8WAw/rGFG2k2QkSwPa735
/VMav7kVA7Uc+X5cIUUsjyxS/p9Ozxbzf/xb5ofM9PxEKeVSUZei/6q5/HIZN3pg
lWLixPp2h7iWbCJ+2v3/c1No56IQpL9PrjgCKOk2sfnUJj32HMdbTIR9vbvbdbWX
8h00EEkEaGbqHl8Suamhqc7JaIvl1qiCZVXuAkrpuzAIBpscm5OrdLtBYYDr0xUH
5d+aUavFPnDoN0c7t0lGRWHmBaH5F98Cl2gh7faeimz5WIdPEIrVNiighTPcm8gQ
f940F6Qf+cC9DXde3TyJRx2rv19HJEbBlU4sl9eMb4O2wgXk8EyU/6JnW7m+vqaT
BF9QYSXyRyrA3UCsvJflK675mkhnnERFCwQ2caajXhPqRgqZp2Mh5qnTqQcImVWB
foqI3+O5tfKcJJINHqc8hQW46nR02Ume3C7i3LlnjOqoAvITepD1A6ZNeUub0Q5i
D14y1Klf+sX6JE5aYS0MCMXkxhkRDuXZSVdAWbLqTgfoantd8eTy/sUpMjzZPzjM
Q9B0o8uU97nK2mAk9KZA/pY7FFUVbM16ljh4aQJYkveNBnjELTRQe0lBCsahYGFg
ZlVS5j6ifTrP4CIdk/hpfbqK8g7wdMyp7MVe8doZ92fr0++yX9nrxSAe7aEKHHtP
mdQ3Hxk7EBN86aTefujbZzRi+nh1QhM0cP0H5HZZycqMzf8EiZGkjzhEnuzAQfCN
eordRkv0d8N1Ni/K6djo+5RUJP61y8LMWQ5FKj/Co9mUhvPpQqvE/XnaJVxfAZix
KG7esz8MPMv9c7VRDcLq40FPexUlgRXjuq4JQAbJzJ9JnDO7RLKXPitOvP4JS4PK
zLk80ZXIxuk+v3TTmsKplQNugPapT1I26OUMGIqI/Fu6SmlQOQrSZndSvC/Gi3xJ
tzPT0g7mFx5b6IRqZhLWZpQn2GyOojMIohXF5fu8qlUUCdtIBX6wUI7FJSxhTDmF
ItNCzwwCISU9EO5EfuK8d9E3pOCfDmj2PhDVHdZNdq6tAMLP/47Mo5xm13hF1Mls
iOEFCYrDzzV6r8IK5nIe/VCz17uIgJM0eVp9OzjVdgl6w0o51TuMuxBgcn/1+Dfy
ztExl9vAbj9LE/LD8/oXfsysURFaqbLJ1OM9aDQ3nn7epK/CILIsYmtGHfc0OGaR
CgBazmgUlpP1ogWZbhVTMz8zAWcHQKtpvfeUee7mH6lR+UBwR5gmJyPfrB9e0KLf
IxXqNSfJiLEGHTydGNyKpWxjZzyG9P5YKjmHF5hRz0fWrxmwfLWizNa6oqgMgx8K
m7ZXMUfynmkrr/oS4U2/DviHRGNbBwrdSsOaI/Xc2+Qtnd5gbrsnJUaHwYprvQhl
sKs0BBfC3S4+lRjbIozg+mpL0NLY2KEWLglJvfY1JPVD5AqlDj8IygU/WfMi/8Kr
6sLgDMBpQTBr4CHobndkmRRJ+BI8trPyiPoU29WDMHg2mlP8Lznuih1uu8lIkKNc
oh1hqJgH/8ET7BO8si7e+pXedyofPKhyZsC3u79LLODl3gpnSEzdxNLrAWAm7Bb4
pWr4bl5/lPFUuQZTwChz6AkEXVEyd+eZI1Y3EOPJbZtyy6qGPRt6+ieFjcMQ29BW
vJIh0I4qC3Oa1aHBt20U/Am+V51SJUuTGu/svzMUmJ7chBnbzxYMKKL5u/qRZ4Fv
5GkoPZe/dJ3R87SbB0siB5H+C7dPkJESosPO/VuiOAE=
`protect END_PROTECTED
