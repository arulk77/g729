`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CzLXqPidC7/gmhvlqitJXGj028Bv92ZTzy4v7OEGsB6p
LmvIHkf4IxoYYi1bsl5fRqCU0PyiMq6FHLDC3j3mbxei8oLAcHxvibKZpGtibrkW
YouLYdxLIPDZ7C48OT2YWe+L2W3ku4awejXNdO34MGuODPWz05bg9WsVDWwFIbRq
Ufu5UEWiBPw7Ru08/Tijf4bYXUflncPFIEudsazcwTZ2oo3Lgl6Ms2CM7UrNTnjm
L9DLl75WJvqeQE5YzKn1nVY+rRtRmP9YuB1OExmg1VRBX/qv+obNcfoqPmkPrnd7
nKa4x3U8wUMWcMleN32XXVVY7VomnP+YyPT3UO27R4ujgtm+gpVyNfKpbXlOJb5b
f85PAzNUOh6apryw+l9mNHEu9+mygkyts65HgkwhBNqT6ICpWIj6iXkT9n1qUFnk
KI+FtiYFwE/o9cSiLAxTuOBSdnj8VWSgzqZRijwXfh0lW20Odc4jdp8NiGbCF890
2qtf787JTFMg+Lk9QSO8UU7tVI+xBJXmnUO21wuJ2OA8cEtstooVkg8WnFJpBK9B
ncqCj1XaUDWQ8mWJH1qdtCivvkjzmKscb+RNa8yAvfpYfxyioNDbY3XeaMCpGOB1
z+k0JI21ZRdwl13yVJhfgDZdwlrHKQSFrneP4GMskxhiqEu/9cOTp/GyFjoKsvKf
ET8MNp3Mtm1907iEWRtb7I9xTFQ05VlfRithVbGXjwdlk8yv6d4/7cMd0iXGWXuJ
ZAerrQeSPnfvaxgChuqaBCiX42vj5EiUX5Ftt3VP+237H3ZMCr/l2nNVHavYbVdq
E5Z4yc4UBV7JoY7Hw/Yh4FBNbSspqGBvYHiRqTOTRjMuccBEMTs2DxZCB+tU4X9n
jR0LFOd+ysLs3SE3OHOkGdBKmGTOUf6cHHyin0tnI7kzTlAcR9+lOPpw2sB9lroE
UeHWcVTQYDKWi9ZZOwICkhTg/lbFVlEj4nITOfQax/1OTLWJ00q3By1F5xEQ4Qus
IPjmdre78/fggW8UyvNZZ8zK7AP/ju/l5Bj16H/81Cs7hReSFKL04odSsc24+TSh
Y1bUtgYl84djdWrNapLE9hcjWwdCoOQM54uKUnZtMuwrLlNUsrFq8gEjRH/Gwt54
8ScKblaBcUFOIX5zT79bk6XOOFjhcq+ZCW+8N7LkZ2/Mb6ryfXimHaYOxyRh3Qx/
4JfeEpQsjLq3R7UA0OoxSDotV/Qq4GgNB/RyvO2byjlvwvGMKDQZfOzgaL6BVgNa
kFFchoXbtsUMLGq3XOwcjoSKCjCiRpi21ryFlDlCpE9VGK8cTSoXmstDRJEKPLfj
tohibzKkJRL2e/0fwKIU7Tew5lZbHOY3iuq+lh0lx6P/mCZr51lEHHeZY09oWNBD
AoEKidIJTtSZt6jtgrycQiPmdoL/5kH5cU/gbediO64=
`protect END_PROTECTED
