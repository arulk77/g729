`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBV264STRRp6Dd4Kim9T7czkUgNT16u4IRenb7gJmkM1
+qHmB7upiQkrn7kgugb8KQm0dqnRvqJ/LqbShzo1LXplUROoyWUV5S3mgOFaTyDS
E5PJ5TOS9S4wcWTn6zwZpw8Oh2jHj5UU0FEiMNouHTrQb+zSWYMwFgIeLgtNcEU1
LdpHBbvIEHXKszLZpUyUIwy9cplkXMS31n6uO/I+lfZoazre6KDudNNQt/WI0v21
CqLOus+hxKD6wnwxqbL2VrFEsuX5hAGnKFzGEzelaYWZrRkuXdi5aX2SqdXe6yKz
10sP9tb8a3tJsTe9QrM+b5WIKcoVqczNaHYWcmeubEI+QbfRvJ8skADDpAX51Vk0
sW+fqgpSPJ+3MDFwjNVp2vdvgFbx7WXaeD+12fklwKAQDUdmb2g5H30TTvj36WQ4
b9t+IrkEMb/8km7IEnGcvCI0BeRnlcDakmNiD39c116Cdp3AJdp+elnCBLhJQ0S2
y8O7wVbZDpPt80mx+EBEWw==
`protect END_PROTECTED
