`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45jRmMO8yr7quvtTun7zXilnUL86Fj/uDX4jHYdTvAWJ
tSX/sjdF/6d57Kj0FhzQJC6AzdvWpjM4DoL34I2xUMbU8LcgWFFZ0hCh37pq0bkE
aNZN8VWBkBdkSsCHFX/9CW7xDdTvwWiI7lRZDP1hoU0nEqlQbF0I7tvqDsDWqbDT
D012F+hHPEqQYyN72Gsc4j0/OMkMsBs2hPWo/OWw6qCRG5qCACxTEioD65bAtRRB
F/PNCTz4ywlPr9RHEITeuLK+XvaRglL+C4EuA4Lt3pQi1GaI2t+Omh0aqnGOGAtG
zO5ysBCdye5hVXFMlTXzMRc0wfWfDP9Ts8RkDbsAuZg7IgAf2Fvwq030nc3+Di7g
SuY4GBfENLVY0Y7VfKYtBiY183yrywz6/aBweb5IHKXuioF1jhtkhDpU34W+cxaK
81oQNu4AS8ChViNNsANnXg==
`protect END_PROTECTED
