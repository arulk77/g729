`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveELEDhj9IhvyajZaHm4zEmWFQw11depqMCJ5gXmVBXpU
c6G7RpxBhJwtecgSUsr6AkdtaAeHCVSMlPHqWPwtdgsffV03je8oF0ynXZiz6TA5
5Uilx80v5KVb0qLd6dh6ifQ4ps2oN0l/Ou8eDjlNzaV12HM14IRS3agrb87Brsbk
c7SQmZqsHghF+uLpmPY+dMaHm51+YJqw86itULxv6QbP1XolIzwCX0k7iWvG/I7P
4uJEi6crk9bkC6xWdx3GG3wPq8h2HX+PPjOlGrJ65J0=
`protect END_PROTECTED
