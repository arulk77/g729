`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLyKLbEIkipX/eeW0hGIMKg0DCcm2rPy5a6fVX156Gk7
wQZ7gwOMrGXOnf8u1Bw0nDlNRgj/3R7ogHGLZgKGeta3fTtkfjTqAleh3LCd40v3
j/G1GxE05EsAghiKBT4usZhNKJZESHwHdrQd9Iz8kH4IySBZkBhF3t/cPFtE8ir8
sYk9rEBCqHr6SLdSj6iXxDe5V9eeWx0BkVxHRfQE2O9Pgxp1oFh7z7n0DbB5bB9V
qB67p4h8kE/W4U7VRuIgdbDT4ndDEYJAXWrEbGpPkcONfS2mAt82domEISDO73Tm
/22Bv1uL5eaP6oSR2MWsKTX6iVsVKUst0Ox9fPV/JBNbCBxHWt2SZ4GGazgILKOH
E0h2JWgR+FH9fquHejK07pyomYD5ocx5DBiLUwCU6d+uJTvRotUBlT40mJOw1IIO
ku5Q9T1fZqN32Oard2Fi9u6Lnxg5MBGNDNmG8jz+xTwL1DPBAnaSIraXJiKWQodk
p67jyzgINfEE9FHqqP7dw5rUYirXeVCzi+87p9dBv1q/5vEt6rnHqcDOQ1U7qWKf
l2OrDYHI/PCAOxD5oF6kaiRXcZ4bscumNX61cADFPzqGH5OSo56KNl75b/Uu2Lh5
eBljkyu0a0ZpADWkF4UxeskflBu3i21N1qv5kG37ceeflhlFMiTF/lRtl04+Agbf
KDLhlibqIgUg0gGvT26jEAnTjQEnW4fa788lty55W6tkqIKHiewAyXc+/G0ZXeyz
VRbLzI7Y8ZJuU7K9N9zHXy3/nBFektpmlZTYG1jTBR9CYI7e9bITtruLnQy1ZPyz
M2u3lrJ/9QJlmvumwXxmX9+vrHmBwFugeTzrHBCTOqsWFk4S8ZNrhsTyfn+DMFQA
CbLwlTwsc7jxHb0uYaEp/i0PaQMXWgCXhiW+nC0t8/5SSi/rsHJFxfHUsutIeNF7
0wrX/n5jQNs5QqpHlXhirAhF0Aw1psJBAuKxVTqxfAQsoRDS5w2Uq5/DJMTLqe3a
9/O/AtH1x7dHG32vYYre9TE4T50rKl0KEfeTQJ+1EbqIw0FXGud4vmIUJf3zLl1f
/JF0YNIT8uCbIF0qeJOdNieScELw4NfQgRoyZzByBPw5PNwu7/dQQmF7VLgIbStW
PIJtjft/C/SpkqlxxnkyMme3sZPjRfleOU+cNBmCALRZFtzfRdLN19qVoejFNzMm
EVSNvcpVYAy+FmLJMSzksfkDEkiD5uNwNr9pa87oHfFUhtO+XqzrjRFkbcmyH8cu
TAGlCUKFtszj2QVcns8MqtkiaV4afwZ6jeHINiTsK+m3TQSlrI8YJZ2WIW3hJDhU
BCZSelMkJPtoGq/Isp1jWW4z++8QtcjRJxHCIpSq6JfEDVkb8BLmgThQwl/T8XiT
MgOnY7m6U2SwY71bqp8+0yOyJqj5Sc5uCJOW+zdcuuysc1PnV4WA701e3p4wHD6b
e5iJDZ+p5fHtolg0XR2u9vzzcjORGz8I/NpAYqhp0XWvz5AgDURTkw5NuizHLEuo
g3M8tr9eIe77tHYrkEw5/PguYI9KX0LZrn9hGGJknUATuIN0VpcCxMIBTNbAkfz6
ohYjdM4b/W353CeeVjnAbQFD54bJifrizRpdql4jTBNa4oWBtHDh+tU+cXEJgPxc
KLjxKZoRAoaTiqHxYsTv8P+oNebBknIZSwDAd2FJDuHueH0H2omg6EBz75lRNmDG
SPpiJhFD4R6sQIEXABqA22o8tWAA4XCdyzXF7U3diyQJYxT4PyH4HQjltIp2fXfx
gMU9x1+cHz34kqiVZcFUqqqT/QCjozmnvP/xMHCHYIj6bna6Oz37zuz5Wesuz+Sy
GBRdIOJHaU7/rNJC0a8i5dSLRlkrf9MjmzmR4K+/ehVoBBRNkemUR5D2iUupbf74
5cQeP/e790TmJ0cXOTjD9V7c9DTEftkUwJKQ/LAiYqYu34xbkOCdlZ7EI5Ziko5E
UwxjykmXU7YX6/telw3+QBl9HqR2wdP7+pBkRyaKFqfc3wYbcqUQExawgY0zrSK+
jj86bxvbLOzUlO02ks+wBcuGJvoaQI71spaU1wa3phQ9RE9//L29Jb15FuWwIWee
nQvrdNdqChUa5oY4sdQpmkY/iG0Uta9yVGuktxdMWAULwFTcJzJ7OnAUFPdrW/yv
Axb2IoF7YfLFlfcN2AmXLO+Bp5P/JYGXrCS+/NulKRrE8dfkP5Tn3bYXg9Bbe/xX
b4kyZDRs9KsXFSnya4LhnFw18UNjmwsmh7LuGnYCN6AqIGDf2Qh3YzsHPwyRhSdj
ZjMjbONsLJ0WfRS0+K9W04l5PTZRXwkrpDqTwEPoMcWCH7co9d0f/Z7gS1SZtOvJ
HZJwOrvJDQfO7GKj4Tq+xIBGuDHQjtBR7WXwUq1so2/FNqNkZS1yneyGz9mOIRT7
OUpHYBNLKfdrnxhWxReWvCJzBAL9uMs0ZQZ+ST+lB8ygO28u95TIdqvrP747Vgd1
Svmi3AF/b1r3qfKLaGA7zsjTknkRmfNeODb9qr+j2b7QOEgZ8G0oh7DwYyKobJyu
wXK45rbJv4F39OKMspXuWPS5M5ZxV42hHFnUJN1eZ/xRb7Th+OVaBag+lgXUsGfe
QV5xprzJ3P827lbsahg91VpGkuhP26W/LjlJI6vrfNoJvpXmSQayiN8+BbRSUrOV
vK8+bEg8lx99YnXDctY+vzJcAeh47cHY67KTxBidCQiJxFFfTBpwlfcAJ+iX8VZL
BoEdKo9yICrUn8OQ+bI5/ylkigRUl/4C9cjgqVeBpzG9FuD4TCk0oCBC/S0fFCIv
CfL6H4IPZJvXmz4DIGCtrz+njChbmoJZkABCqbz1NttPKROcg8teNilM95ayvpQo
DBErrfYxFsLLEuEyFxKC87k3woyFVNezTMfNnQr6v7yg7l96NQUAv7JThlS7c4O7
QALlIs/Mt8lAQCy1zsBAJfp/ziedLvMLD3jWwI2xZdvdz1yKIy8GmkJqsXowI+VG
7AdBukrDO0h0yeaYcLRetGBQ44TpOaZuw9Ap4SSA+eLwL9hCY3u22fgzLk92WswB
Z0Q4P/dtgfd7wNE5aBWzb0H7Vz9/CuVQwr6oUZ40Fm/W1v0cYrbnclVvWtMW/tp0
lyVv3Y62OAV39+C5f4dnAQx3dehHjsUy7ZkZ3gtOMh52VN7MpSZ6/NPyC+EPyb4U
OZW9GLZCjqxB4CnA/vYRf6/KuWaP36yNKfxhPXMobdnkbAAPWdJmtHaiqEeO8IHM
PFd0+MAV1sdeouNvSBYt0Y6sTkMAE3p04ihuDxmJhMo2wexXjleALr39nK5LZn1D
oum61b0eCS9NwfFhszVtgXhvj5B21YyYN4amb04gbBJGF0zdBvmRjbtRE5S2zUFI
gNmEwVudqTuhnIN+rGNVWK1mknU5asUCt2il39j4nYDNSNdPQyyyJrPpzUk335hv
pC9JP66KPtE6Kj/opvgZ1wo308QhLbykQQcRPd0LlwILbWXJo5HPR+wWpPLFSSa1
SXb1to2ZDObPFbfOM2fAA1di/ruKd9lR3KQDcz843ikJ7ei8krGq1Fe/yadkRbc3
uxpUSGN6DeHi6arcoggIgrIzmHJWnM6XkAPEbUBjHhwQye91DltlAsZTrOOUKt9+
4oBzwqHFxvGz7s+whAKyFF0zn5CJfdwzJNxdUzjrdJ4d8+0krDzEUoPQldx1/b9i
x85TaRiBgqel6Uuaxe9kAr3l3QtXfU5ftTu0vmkH1YcQVgORbaaySrexXSt/6EMc
tbo6m+3hAdBHg2/t+FMlcQ2V72aKu+CwXmaYQldyxr+PpUueUkvJL+wrOKB0Y/VL
7s+qLfNN0afhwor6mHCFe5KCDLlQQEO/ABMQpHv+FQ/jj+u73p8zT/1+y7XT2+Ux
7I+SIwTuM5MwJd/wKy9udBWOJJgf1Qk13K1aPcYCsf1P4Uc/K9vomWVT5wm9lnMy
zEieHVVoie8bNTGs9eqeNpyCfcfbKBOPKwcMxzal1TkYXfj4oW/3CZOCFlPwYDmt
Tzqts0w+Io7eS7+dCcO9d9sKFBUB9Dk3D3aaXLy8pPrHB3iDzErFRrN3sQWAstYq
su4zqpxsMnmOF7shC3ace9clY8hfNkagWKBS3b8iwS0n+fWGsF7dvQW1RWXqAzXH
1GSXM7qNwsk40FIooe3ttu0k5PB9dgENj/JNk2wHrZqZ70Y9pACdYK7VIMfYnvnC
QA6p8YjvqG7gNJb4jup1pck4RofdI34u7rjeJYw3+GI6FYlpGxPKpmC5Vw29jSfs
F2A5mIxSrMecRG+D4E5XvByydSguJI228cdi3kIKV6+/4JZxrsT/wncOF+YXFq1N
Ckk7bYkRE/Pzefr9GeMSTvuhxUDrtyKKC5A58gIaWrOBe8WOzhA/Hgw05eyBEJiU
yx2nN123xM7FnwXCwlxgCkzoKVc1g2ljjjpNy4ghb4XQreh7cabWwuhlMgMfFnkF
62QUiqQvFGuceFkd0PSBV5jsprzPnOnSUFP1RAEk9YewLub1WXwRuWyER3qzzJvz
HM0xCk4u09rL+35RXixMzveHV3LQ4Gvf0xrYR11FcPxx9fok4DL5hT3GMwOVHcdU
MrmuQDhCy+Boo/qwH+qP3E3aOmZmJMr+drlwnQVqKxM/tZI2xS565N9yQhMIvfXr
xeg3uSS0kdPNxCGCk9AAs6HsLlGZ0vqbE8/wQT0fOrIjJAogjQGECE4jTuLUggk5
kEI05p0hXwanUZOfaH6cXOPCxzzNKDMjmEsJNHEUI7sFZoqdPXNwmkj9IOv5Nw/I
/vla3Y8DLRLSdG76rlou8vUu/EgF6LzEuHiLk/4xcKnayR5dfOGb8XPN8I+HTxrP
`protect END_PROTECTED
