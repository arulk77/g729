`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aYf364kDYmq5V0I+MQXb+VKpRJa0Ze6J+YGsxcFB4U0N
tnKEFp480nTzY7l+cJ7HbKdxKGS2MpAnpZBAiWd42AWO435dsOPMsATWzl+bNchS
PWHZflUrVOHG4QXUbCl7JVxZW+bw89WkW2brJ3yGGY8W6Wt1YB0Y4AWqdeWn2atT
IMf6IwOe7T/HNBGBwAmK4ddrKayoBF3d9v1Svx5Mug8/DwlGzHz0XfPjH5QxhR+6
GWV6DKekh5Zxe2PxYEKZ/mohE0Il5n2Xqqp7mQeEt4ufuuAsbDyAu3740nwoCqAI
Uypb2oRdp7aiiDHGmBdRuwGwAjrpJkd44eqNh3gAnUB28N7fgIv4QfPoKJojcMn+
tU9eiHMS1+WDDpJBpDJHrG63ir61dgNgn60UQVSY1ZOkoI6QhvmxKKpbLI4Aqh9G
8OZF2XULpTK5m96x1vExkF1dATckF8Xki1odW+35BF/TTjE/16ccTTZzm7AkvRVI
M+0DRP5MZzSX2Uax+yOsvSZCGhMsfL6bVPg/qccJdJs=
`protect END_PROTECTED
