`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
83wvwHJHdOW6+Q/6dJfBK5oG+S6N5WsUtlLQF4YP2TJBv92d+4Pz2FyP73vnMeRU
0Go4UGY6NSK/u8barjhj8J1IpJdFjO2wThBmrVihYcseQkGOemhYunD4Lios/KY2
igKmCk0A+3ckMS6m447pVCjXuMWcFRevNU8AzDhPUeZp1hpoNna6K6a5JDC3lhcM
tWk5Ra9yZSMoJJssUp1KbHd1N4FYW69P+pKmfDIqaxs=
`protect END_PROTECTED
