`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSB5zORaO0kAI6TBt456HXVpC5N4sY95iIbdK6+XEY9t
Cpyo0vfaiC8tDLbdU0wdpERPIGjTfnsVIuOgWAZcBr16Iw46bmiVzUzW3hIxNLfG
thqUFPextmvTzy3w2YsP98paaUtwp/KC825wXGncupHTYscD2DCT5cNsdfBnd+BL
o00eH3ArwNDOr500oOWmZn0GhFztFu7pExlz38P1Ge6S4/LxBbWiBibdw1JCSv8S
Z0vJzveJ19+ZWKfTZieTsX7i7yjAFzsuh1wtzTJ93/BaXO1+iA3CXvY/1WorSAqv
BZVB8WCU5OZLIO1jKKwJV1LDYT+NbciTiq4PMEmI7TzSrt7y0Wz0YnElDz5TkP+g
bffNcmEfNgqhO8XtpHSaAOpEZAhee0mxkxN0XFUuzkuagbvJtIPvxVa5rKJCvQ4v
PO/C27Upa9CPZ1gKnUVNS1wAWz7zJFd2bWRCzv1RYMRmTrA4PjxXT6YCm7e21ebH
fWtBb9tCEbo5cUkNc2wLsmDSh3xLmXSbMkVEOSB9JxVsLWjOt/JAm45DlC2Gq3Zc
hAKOcriiAlqMhuzYAE5G9v6qDU8rHMX4RrDX0S3ZEe281AKTjddUhb3mGbSvrChG
KiVLKjr1DxgiU9exLVUfRnTonspftv5V4JwMkgDaOdwF7EazCsMr/3xpSRVyhUYt
n1jQKnIoTgJbO2fr7vDiegwz4RjivYDCN7W2xoqB8/y7wNT+NiDQQ8fZwE6Zpxe/
57ubTIyEPOOMqaB81gGOcRWeZxa0/KdSON6jzvNhSLKXBveZmbkFMSau+HahHvsI
mOowhlYaFpwGTaomnNwpF3hVbMCbh4ohkRe/XOrlLPzx7FFptEVKZ9eUUQn4tNHy
5G/TMJ+Jj0fgrzO07hRVrt3zjmWrpyPAOtMcqH+wOHLIMRzC3FfWCqktpEIv9d/n
yvRbvMaBYZ3Vo3tK81G4PkirbTIttsJusqPuI8ALp79ZT7LFU4Fs0p53mKaIrSeP
gMPIBDaBOBzDmp8FvUYm64qmMEWsrU7FDxQWghjYK/YiTp2GZURMWzLw3AwaDh8p
c+vd4sh1yv5+g/63Nf3m9qdRPqmQU1O76UInVGmApOqB53hw7I4H5qUnnIeTqzdc
BCYHcobsrslyQS5I8osmth63xoPW6fi2su4iEPDoas7vXKFlbTWc3muVepWmzCZW
iXPvG2jd57tyOMuj4AHzaXSJAatQpxmuwef0iqja7rGVPjmQpC0Gsgd4gfZThyND
ApGacnqpCBrYnwzUc7Vi4yHoxmmgXKlvUnkj8nxLNc7ZLjpuHrvWmEzZ4VCpqXO0
1tt2OxR6aiyeeWSNdzLxOWRfIJBq0Z1YmKTmb9leSz/TTyZ5oFuOkDjnnbAms8mR
ycmey9DcgBfOabaHh0gDw/dG1YPm7Rfe67JoGpa08f3UUYbxg39qCqZqMrF3b7gK
pM+VABm28Z/lYZ789lOPrc/Czu4xNtsT2uz5uAI7g2/CQQgncjBE9xWc7okDynwQ
5VK0sDRqWmlyASptfePyDkV5cRM8ZFmCVmr2Py9cv/50zP3EiTksw/L83A0QLCSP
0X/xNGrRD1j6Vw/5kx+jqUjJLpnYuVyyj8K72co3e2qNnXwPIcT8MZPWjhRZRGsN
2S44fQ0sUoM4WMWUJ78CfFx1Tmc3C0uNXOvCCGtTNKqJBb6uiTXpb0SvooMdGkiL
RXzNdf4SUaGPJ++MsruHwEF1MsaeX6JBG4U+sPYfIXaGbP/6+B039moSXKnXx55c
r7KfL2OvoTn2lJz9uM9bOPPeYcHqK2d0T8VmgzYt+zS+/HASfRRPPZaLo6ZAZnXw
uImKWw8LVklaral33lWhl6JPqKzHAToHMmNdmqTrtMdmSIMd1nsnAtNE6vJrEhQM
RJoKy8QAWUlHwcJ+zwQxcQhOXsKnW9bixECXXkIjikdaKAAbDKsIXC+Ed/4TqbMT
`protect END_PROTECTED
