`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4dm4AHastDqRBFj6Fz41cm4deICy1SZOLzKWHGMAgB0cq
9rcCD84G6noh0UkKUD8hsfjWFLaXkfCH/xJdaK5fY56wcaFOwhMPfuh40mOU45vm
5O9tNFpey2FK81s0SfqDOnXNmho772179kNKoDkI2yV7S/tDutGOmAszavAXWRJU
QkbZJ8g1vLad3V4YGF6v3XjNwC4NJ87FlJ/oJSgCWrJaeqzuv9lx24coOz61HoWM
V/7I8cpFt6QEzMI74dDMFaHoI8sHIO+tT0/WLDhAkswdLUxRBsmvoWW2dAZCSPf/
`protect END_PROTECTED
