`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDARV3mnor7P//yVlll9rb3yDdOcOxI1oe3YHw/V+BEZUV
Urcn5orpmODXeDg9K40o19DY8629naxzFrTVSR8YNBbZfq+lPoV+ZsHDShqT5t8R
/bakHljFrYP5HOYFgjrblek8LXfYGHhiQawM5/dSCL3BJlMwnh/ZyUnGZCFcfn/Y
1Q9mkdoW+cDsQ8xmEoWYsRpSPeqeIG/RCYj3UXM8z6c6M7A3J/5YE1w6fqHAsNzS
K2YrDqec7OxLVyO+8fgTjoTs5mtUpnl/PTSyuH3y8MHJUKZ4npT7PqAkYqiO8Vrt
iLjfvQz/YVROfd0GGIneOKzRcfJNhB4+oJcPRK7xsASIDCVe5Tqsr2eNYGiafC+h
q8OxPL6RBsM9X46KwRjEaWzA43ctEZbbur873F3IlSLzbEHKL/01sB3LbnKo+ZN+
W5a6J7BBCfdwrOklqBmGft/2NHXEUU66gvgbuQqbc8n6KHe+LpqlOJXwAzt+gIO3
9C8dCdNZeQa9cBZzwhdeXwqb0IWfWI4HRkbb6EwUqmQFpgJOxeq5ZyCJ6i7GsvPG
0xD2rxB46UZ/CWHFSgRxkf0Q4vA0pK1BlISGTw9OC2IGnRT24TKTHyBJNiykOcd/
FiLspR8CiTxdG4LEQeCuOJ5TJlV6+13PeoNtYVdOuEjzU5lSSvonTIzzJerv4k1z
ASJ8o7ksWukYPuWlIU0gfaF7SwePydaCmIzZ9ZLqAG+QZHOtkHvvDoG8pdOHrUHD
bScHnnAfuqUxHFgEIrQwyDRYRDpteOOmtIPhRHKRJiYWsAkXzXZatn51KpuPjF8V
IEBNNmca68nu5IiFnJJFjjS8VbEdJtqWRGBL/7YJYZmWXQgbxcTqncwU7OtUUlz9
lqcZuYhUh1dEAOpFA7wEv3zguFdQjDcSuwrbmi0b82ZZE1k2BY4SwGl6Va3r64qZ
vrhb/gYKkFBaN0Z3TxXXF+5yPLBLAkBMGjlBkpxZdGW/EItl1sZ7W+bh6Rq2RgWm
JZb3PcvfULDhM09iPXQEzdEDt7OAtiybtsv6165BJ/IPT9GWMExZYaINiebkVjex
pTWIwmSSBENWU/VS0Y84D+LnoZg9nfpw3nyxbw2NllNwyI/jzDybzWIm8wb70p1h
TEBGanHVzA+7NjBN4otmp5tZhz6pe+G3Ed2AUch/O2HyFF0LHLG6bUSZhd8PIW9V
vtFLJJEZphSp//eZJVBrcyYAX78QLhzkTcXy85wf1NrmlbNSSWbFSLZAJUdJrQDg
wm/9guEl12nhXmJAw/GWMIbn/oagmA68rGBEa+jnTlkpj3RzWPWlkVIWO8pdVq6+
MMQhOShISbRknHYVPim0QDW83o7j6vkz0gpGBT3y36fplKyeBQvSw54L3gQ/m6j1
k5M9za6sPrELy4hKk3pKAeZbdgLIfpy2PC6DoLV9byBnIXls5NQUwRqBUY57UueM
BxW2n17yE53+dtk5rsABmXqV1P8+pn6jTYSR8iFOMChCy2wwAIG1pTCNhz+QU7k6
X0OKsKz5CMIvMOJARCEOcUB65gZHcI2XdZfF+5HTqwxJHCJdsCX/NF8kWoUS0EI0
qE0SpFMkjpAboiBKALZXwjtdrU9oPP7zH3r5V+mTOVM3LHzsBewoQF50eLJ8H6wL
WsaFEoHaRgvi/q7th7ici/vNC1GyuOljrPVaFf448+MjblET6r7W+DRvKkwtllu1
FVvV5iKTxmCRuFUpBJPXWf7ARDu30RtZpX3fEodQrs243Xx2E+M6Nsh/h3A+fMzx
6EOLQJPHgSmGl/VAWy6gSZEWaPtYVPHkBMFGRAFp4INMMdcsKi+OG3wkNHn82/kp
6L/KPLsH7+5ctIeBFr+4a0X3kiQM5ILLdZeuf6olZIUPa/uBqIbGjPHkk3W5L2GS
TKljyO49XYDiNsMBWBEeYgde2oQOI46qPk0XHHaRGdoSGCXgedxDBNua9bbzy7RH
P+4KeSnj5IEOQd87/GGfYg+3B0rur6UIls0aJ32BTgKhBUo3Dlv2yeuIHpYkoW0C
VJHwm1RJUgq9MBZjfV1HPaZtNxWd2R0BvQtzgYc/lVLIEn/AZ69H59PBiTExi3PS
l2d8qIfkqj22Y3rw58pVAckWcLswlLKcHfBKvwmggwzf2/xiMcT3Oyox2C8b8zN/
21qid/f9Xahu7qf/TUI1cqZrzbXlMsMurs4u0YHzsgpQsbT1iZfXWiSIiC1lsMrM
fphBjmcFxB7Un5ghyYYYjS5bhq/gnHTVwVADX270cvA0yR/seyZ0j/NkRnSMvU8r
GHyLR7eGjzsliSCKAkxY97IloZ8ceDicW/YcwA4I7O4qH9rbSDKUN8zx9rPZfvnW
exqw+KKOAoYwkyEbh9ggc+LLF3V1VW1b/MP3DAgMM56FCy9ZKF7pQwFLKIxPo/sY
vqIXyX2PjAvvQaQ4SYkSEyEYXsMh0DXgh/XaWvii4CuugAKNGSpSdazawxVJIwXa
p2RMNxtDdVV2oXBLAItHtClN8A5ywzvdVLXg4xYDqmyccTgo4K0+5Uk5xQAzzcXY
g7pXwq+ZIBUN9V8DCy+U+a8Aw+z2fC++rVHklWyGrCsI35pvtSG7IsdSK3aT2OUu
kbmNQ9f9Ozd5mJIx8WWKupE5HMlCuo9dBPvuyFTMLlBirVowNjKKiXgROjHvkkpJ
QkRjHO4+Y1UCxeU/6JGRWwR7Zp4z8pf+7fPLdm7Gdvxkzhxj85ttc8uJWdBOL7BD
cdd/1qXvZMl3wj0Bhs8qJ8MgnXdbyTS0it1gMkfVtDPtvVWlnwn6RoCKvXrQGuyx
`protect END_PROTECTED
