`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jkR4h6TZdnrSHPa1WPizYK9MrJoYFeQ8lystsXR5++VI7Amn+XwP4Y6R8UHXVEMX
0Y5vXtaqMnZ/C2TkJ5bZkD1bX2t9eJWUO6LgIZWnuSbnJX70E3T0qefMEmcrGgOF
WFMiYNHEnm8lhy2xLLytopCQQWZiUaV8s96e0gL64LLicNcU+0im9SrBht6ywqlp
LVUcFV/cMglXy25NKbzgEzXIsD0GgLdME0z7EyYpEOC0+Mu8iQtDDyjIa8cE/h6f
fqerEc8Cod0LGFW1Y2VcefXekbs95dU7qiZmokaDE0lCeYEYdPk+tjCy22q1iWRJ
53tmOSFalAHtJidmASVhhXIjsKFieR+sXTQDHeUK1mLpeixr51NzuvI10j8skYhk
22kYEHVXHkFERgiYYguVO+xkbaR+84FNeqA9MetwlL0=
`protect END_PROTECTED
