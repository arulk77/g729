`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mzvg7cXykaGwoxwMN1M23oncO9ZGCCxY3QbcABI+yuY0mSV0LytpMdKYM49niUW7
QiZREXsXaTZMkwnBHnNTfX/2nUpZX5/wBq+Qe0MXDIxDGxee3ewEeJeg3GHewyTL
0Q5+DYS2icRol9zoqG8P0k06FUEFkOA8U8/td3FWyC3pSNY7LTscfHcEKPWi5to9
+JNlgOayGHWdlKvpAryMfi3b9w+zhLzYlSq9nP5001f7BqrTKGWgKW7hqyvMNZXD
1IDVyQMrG9YNJhhf/OBxBmYz+PSfm4k1rPw8YJIXZsXik49IToqZ4cyNTr3W3ITG
HFg8xIhNDTwaps6n9+uyz4CT74h4G0E3Gipw5M3Zr6zv+mi/MQYVyIIF+fYiKN9q
o8Q16n+BOla/iEDKFk7bDjpyWJyu9s3SVmrH2tckwGOTmKO1WWFRwxx26LiFZIrt
8zM//OCx+t1D09zrMu5KtybRKanFl5GzIE609yUSkqja8GH3tVZ5TuTrr7Jo0tDd
ZV7Sir07vrWPZR44DLtC7XM4BJw3Xhv1AjQqw1qHlpRBsLUK0JNyXIvGyFQu5Vwp
1ovZojzPbdGyIK0ySZf6VQQTvFM122G/l8yK9L9YW29SyE2cC4rHO5VzoeKCT5kn
VfZVqQu2H3YrVwEKZwp79rhUdCKx8ACi81NxBmJXpC8aq4yA3fOQRx27Dg1O8QKF
hr6ND261yo610cvIyN/pCeTgoQNgTuziM8lsVEoh4jgUj0pUBKHQhusiXcUXtJib
ITom8WNXFJ7nrfR37z6Zlflo8hlAMm9ZFEAmRF9VfVvpesuaMcDSRc4p6m8V63iw
FKFMzq/VXQh+RwdKjXLNckuamuzegHWLNoTmj4w+RmoyCStdGC7hEpN0tV0dXnD8
WepMp0gLthaS1kCR2ImLb5EIT6nvuAitzm1svz6jiIln6peafAFwoPdg1q8OUl0V
AvP0VA5KCwtDDCmddct/PP0MagugcuN5FZ9HdRBpe21CVqSGsiR2qGca+kC+bjqi
wUAQx1RyLAIpOf9t6Ye8trsvPaw/ja8cvvZr62T7cBoAnoo/PPtApWW7atWDPrw4
7H7Q3l9jBU6+Uw23AfqmXkfhedZm3d6qJOu7zO/0BZvonAAObbpGoEQmIdwRWHCr
0z/DbWtrSH82b4qplqC6cgMi0Krltxb9ue+25m0OgDEaueXh/l7J5mVn5n1+4Cdk
9VF+Aydl7U55sxdK9QmucFi7ilI2Dsk98Y+Yj9glHooQjobnTr0F8fAlp64AjFsc
11+PE0+AsWg3BpdxCYxM+LXg/ShrZpU1pP55lkCqC579kfSqecXrslM48DKL1u2t
KWNcfZ0Tbtob1xJiI/PyO2d+p0jBfLppCH4C2g+jecdKutpbnbRT1dgCBqgSI+8Y
2g2hWoD6FbLQ1rXlByXBOy+yH9anEf/snTaUu64bk3uWko8T9jf9uU+j27I/bMN4
dT43THT87Cchr0M1tlhiVdY0axOn6BHsjERQOgQwkZwQpGkyK4sMdIifh3S/cywo
YnSWFlCuGwcCAEr/yKTE2JwOe0+qz9Q66d+UH5BPZwflUV4AV4HRrcuYyfju8HPu
q6k+dq5o76bRmsa/DpY8nlpZ0qZexwxur7cjTyfze/KOpioPcBQPzjFlpfHdbhvn
s0Y3DhGyUYYFdJ1t4ggmMW/VLCiy3Pr6OUR1F3CaAYzSzCM6RVUmtlUFmIMOBrd7
qYK5nkUwWizkh/o9Rl9g2w8EzbGBI4zeJiQjJtl7VTq/R2LqZP7pNv5a0bD/odKg
rGcbXMH6svZ+aCc7uzfrNGLrStTR3svDf2L/FW5L2nTjQv9cFcGX5eUa7dC+0NOn
NkHM3tgIyVnQDboerQkJJVJtokcOKvBdFQ6VxWtU1gm0fVGLKOHmTrxWSOsyHMlf
/C7zp5ONhZFQmdyChwYZeNtbSDM0JsbXU4/ysB/V/bSWMe7lwFZw0qiQZjxqMQUS
rf+XxP+dWm1VH4TLkiQTiegiWRG6cWlfQfdbDShmU5l6Wldp5G0h10Syq3oTp90J
Gw9NS4mtTNC6/qa1zHbjVvwb/CP4w7ZIfkQinZkl4UdYbkYbXOdIASVxkYwNKPQs
fuObSHBiRdD73hmRI3llNq7UkOEfhj3QY3sfWvzg3wf6VT2MWOIdW9inz/7ftDc3
1xwl3sGUCtOb8XbiwVzRbS6DQYKrQVpkajV45iFY+XKFstleIT+8bdm6J9sfrT7q
9g/ewUy8GunYP9mgTyC+3a1aJuqcj2xyHcuVT6F9J+I/tD75vor8sUOes3EOSC/V
6fUA6ausiYwxCMehEz/gd0Tj9WmXLIctCZrU5ZBZzbIfpSKRU28DvZhV0ap9b3L+
MoNHNJ7Wd0LyTFgcGCI0UaSgXT0SeC5g8PIYzB+Jj0jKV+F3OCAdBRAzJ/04O9IV
9QUj8TPi3jiSIfSNl1K717R7oh6N/RZ0kJdU++n5r36a+XL6PlnIbHtg+TO19lm6
1rMSJvZuVYqRp69YrOmr+AaI4A40HJg43xWDj5ARIlWxuRrGUxEg3pMGbvFauwng
yiPOM3z1GeY9XMUONcc4Ltxvu+NbBTJZFGzU0twtf0Zvbg90jl9LEoB2vMoiDfs+
cNaOa/1kM9fhBjBmS9pHKABwOeEuaMxTk3bMRMATzckHyNGrWE71zYvfnRoktsSz
fK5DMdItzQ9sKYfvngUetTe7pz4cn/lR4HcAJjenCxsw/Fh9/JgC6xpR0dsAB7ks
AHwgfxWYTkJehn/bn1P9wq0RTTq5AC/9mDgjioEGAOk3v//52Kw98IwBpd9TUXjf
CIa4ODghZzTS5ViFHgEJgNOh4AF8nxWU/UC3k/4wjIDAL8KLiv5o3SihmzdvBGrv
+IDPedh9zKa/h4OySnzjPNx4e9Q5lFPi1ShRLS1t15D0eRfIsgJhVNgX+jZeVyJd
IPLciTzp9e6vPWJ52dXNbp/7qpVOUkvCTMzkY61jBSDHjDOzYqB4g/sDw0zhkJq8
TU0Zixgt92oHrYIty1FSdqgMB3dhq9myiqtg38MRP4gRp71S3KVIlu8Hx5W9MqcG
DvrXmsNNqVsZNfJIdxfu+Wvi0lCUE/AOsk/L/xYLlzbCoYXaEOaX9lX4N8g2/R//
EPIw285v7kTtmFojw8Kody4q2XeUGCaDeWR+SE6USEmMuPMwYlrnA3iiIqGlPqdJ
iKDQsHfKY4wOVVD3G5AhUdE77xX3rHeRLypPEYSTtDsiTFcMeuhonn+ni4VgMbQ5
QpXU7MFuD4CCO7+sP/b/HwMJYh9voBwju8rtyDt+akNSX6MnBDgsI3I5Gh/EYbyx
o/l4ULF1rBOCpQogIDLcrcJX9o40rhDgUqFZWTZ/qoC6viYoC/ziYs6XUqYCXKCc
J+pAP8T8O8EFhWt4XHziKn+HSWZXAITfY98akjJgX4Y6+64eUL8N0rhfJhv5gXLF
wsuIFwd9R3cVyBmaovD7vr6dvqdv2oUS1eYX8xCwt7JcOfUlk6zZ0scn6YWUiyc0
h9BG1A8C1lp+NGsyfobY7MONWxA+mKg7ZyZb9ItvV3HbXLOrzvJSKu86BmMejE2f
fpUZ/z6KJv5JnkXaUxs0wN3B8sEj7QgIJTqFKWJ7GIrzskgIHrMqLRKNEWbi2exy
+S8F8eJN4BaeKjAVrG/WY9GZYGb9hUOmZGrvRoB+ZU9gaAsJ8xPO3eVe2icF25rg
FHVX/o8eC3nhOVggcYPIo/sq5zT1mhvoghgVmHgMAgIU4gKQO6J9oBFrF7uMlpTZ
3kSSBa8r/3FaFwBkIs5no+I6kznWk2qrh75OFbu+weNpCujQY+NDdy3dMXAAm8rY
cERLMP54Wix0welSYgzyy6gg7TKZlwUANrYrkLBeMrjjiGtKApMmVL02zy/r+hQb
NdVJuClUgl1nrT2f3XkD5ujpGeR/7p5THwFwlYLd3IUhN9SbbvAoux0G+Ro01xgB
Mk/yGTQsVpIiDFPG9wCCikRi2S36WkftySnj1arEtrD6gBSOsnFPdwqZNwnD2jFp
lfgV9nspYbW80EMPdQgBiPRHbrZuGzem5Tl693Is+YYocJ+etgySxzX9lvGceiUn
56nslKeFR25uIkInWBMhAvZ2j/e6/vxvOchH8w03g2l+ggMDtQOp0qmBqOQZXAdZ
iMaSMVGptlFGmFlHYq0UE1KDyYiopdwgsOJsQ2BxiLKnj9/WAiyfxX/X+BMX+gt/
QkefhQTefk0fyymPYbgFRRQzR06zi5v+vSv/wnhCmW1HBvwIpwzrRrhJTe75Df+b
cwIVQykKmNCEAmtTV3GDPs5rALqNyLaBc69/ZvN5CqX3SLE/fdL/fCQhlKVfAkiy
BvXhe//u8Bd6s4K2Te3M5fXqPya//peZlogKJL/SyN/YX1p8JIFVwkGPCp57xILh
6VyjHfegstI6EJQpNGk4CUAmPbYEF6a0OsRrxp4bND1TnE93YGPTvLl/LMZbIXkR
34CKsCR/ZExj5GFkP7sI5V0p+sgRRIsRIhbHwvLtj/nQZtbFFMJFsTjmFkFS5CVg
RUKTsboC74gvKd59RV7BNrC+AgwCrdqtSW7g63ErxCZ++wFR7JtMSN6YSNaN92wY
rR7ehe8mNfGPpwIOIi8O9vkrlapOoDKryh8SqOOQyIyuF4xMowrA1JSc2+bOeav6
XzTK3Q4Hl7rmnVbMI8Lu5QtCizPOjcXW61TIs2XkA+Y3kRbNv/u/cQeLvDyailRv
F3i5PLY+WeCt7iKjL2xwWLy7wSMj4aY+5WDXzni/Xcd8/cCOjjc7FTFhbF6ut5V7
MFtiYnhIR3VBo0NDZq25eWKh4hIqKDhXOFxFR5it9q8gZEA9iNYcSqMZiTxIknjJ
br4nPUXOjttuRvSVVBQmB8i7rO4quCHnCMWTESbyxst3rm1g1oZay0ZIYukNTkt7
ionNONE9PCnIGJD43m0mIoqmc8HCRC6ggLA/HruaLM523s36lVRTrjQWVXE2OMRn
c6j8Fq7Vs2S7tFpBruW0hcrocmdW8NKWpITD1urUpi45erxigPW7NW0ljAcFj6mi
pVKNW3xrTN/jUX3QB+7Mp1BWLpnaBLZNADXP6pIHMfHvBsoofqRgzSyH8FD1y48o
iGn+EeqAW90/J3VYp4iw/cjuUgbYeS9XHlBkiaLVu3qyT1Eto4Zu5JqvMVx7HwSx
H4vKCzjqaYJ4zF7YyQ9CNkMA8QSvt3weKbX+un4vWD5adLF0Jf/CA62JRKy046NP
8bm6X0yxVNdYd8Yx9Re3Dr2Kmnvgh53CWQzuBCXsR0zcVH3vcsw5vO5SBWMbM8hR
TyFfRTT0TKMKkG4L1khFXiVDwMvSITcPLZrl2+nSHrko7BRz7ePYx0YwGV0TA1s5
Yr106KQhp5H8u0hIS7kgm+LZEIUS4zARIDgXQnbhuonOwXhKEMxh58kp0RlQsYih
yBW2wuqGU7b/J4CvI/DWuO78qMjocDwSCuTG7UxJzA/1EqiwBJHAYqoM8ysSV5XT
Y+qmY9+4xezezBRPXQTzFx7J7Dw5GF2AZP6yTNObItb/J9eRu6ajysRLWuRxKPaK
YizvgfcxTZ1GRPY78OjKWMZgsWvHM/KghXJwJpYDi6N45Syp60vTSof3dWIAm1lO
1ixRDlynsNVh98L1mXAFYlvrddn6Slk+8VZBMz3SmJJ33ns71TiTQ4oLM90K6BL/
oF9a/5X6EuNGt2ddNrTKTdidIbFTmEd8AmiwFrzwl/eybA7i2o3Im0QEU+lQ6BVF
`protect END_PROTECTED
