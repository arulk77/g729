`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pjEWniVDnMDKO30v1x5SaUeMNwDYBbgSGM1DD+P5iqQy/KfiotoxL0cKqA5ovP3x
Hnx+vu3u4fMhNQo41vo0qDxG3Cw5nqNoCukCvjyqF5cKQKOZcl8jq3o2zBQJe6OS
eYW7GUDmUilrD/aHL/wWOaRotV75M9vaHw7HfMlU994jH8mHs/QEjnj+oDaj6XtJ
CLAqzyVoVhcUBOqgJhOjwlorqoqCDdyemZHAivmz+NrEz+pdr90GTWCa10pc2Db/
HML8wZAso7AVxPiMSXvYr3eybHyHP81iwmap41VsDjR8ZjwsIJXzB0S1QtBTHL5D
XPU4VW5bKUl0ii8/vbNoKbmLb+Ev3w2PAMMLX2MoBsg=
`protect END_PROTECTED
