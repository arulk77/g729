`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
b4/LScsb+PdHhclb5UIsFaokGOTN7d1u4XDhwv1K/tVKrCjxJxBCdktuRO5Mf2uy
RU19wCKqq2X0+IpIUzKcv+BtoWHFlzUnydfwt180Ekk5UsD86jmPbq8d9csSSs2/
yypuHkTln+km/IYcFVPVkysUKwsP4L2KfymQkL+0pU/p9Drs6o/JzMvlyW8+9r1f
`protect END_PROTECTED
