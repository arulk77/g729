`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHoLqjrjfLdLNi3t1gEW9PlCyS1h01esO99PfpkyLJ3Q
DoPUPiD6EbqbAIhlBfDvKYMsTm89pYC6ZeUFctNQp8mQmYwxLtW7ypMRkDdF4GEG
oQ5+vzy6l1iqFzm9c85QiUjnDLB9FDRxy3rUiGJByiIjKpj6h7H9PiNyWuE9e9ga
lQqCOZD1X4I8GbbZIqXpoA==
`protect END_PROTECTED
