`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xyvuHe6eJODWysAF8Qe99xQWzRwetdU3rwsYZcftkXx
Ic1r5gciOVRvL1JpYDSwpd6L3jhK/sv+952DaXowGYtXuz3w+sjpxhwF3McROW8q
ia0gv0YqePzOmenRrTFvZXW9cFHNOSCJHvMyWmlg/NQ6yxdN8uzEPm+XvuWOSxHn
InohfRinA/ozfh+irFCO8UiQicLUGaBDS2l8XUIm2TewA8F8BWDRuTYXQfK4lPev
JGPVXwa552Hdh8Td27yn9al8jqWzR4WGb9o+ouE2jUSuRMMaLN5/w+++LGxfe5ZL
dlG/FS1sFD+nHqEhwQ2NSQ==
`protect END_PROTECTED
