`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcOHWiJofcvC2R8wVU7I3pcBRJN6obgMGFRxWO6/I9mqw
5xsKCTc9Ed385cN07/fSQcYfYBE/+h+0uQ3E80zUIawOCTmkv8ChMDd30mAfv874
gkaU2aqzp0XkwCyhY1izLA8YkjQymEgg3tqVdTPhZFx/GHWt8xJNkiBHJ8S5DWwa
E0HjlDQ2eMLeYATzC2SMLd/HwuaBdeykP4vW4jqRPD1I0S/BNlpzZlq1ZcMJdmM3
kr7al9CKYOD4Vm6IVpDmNCt9C0qxYqOHcdjj6DTM8s9125qSVxgjX6l/yAS5BkHa
9Opy0Nn5eQN0Aw9Kv0Wn/d9VZItkP5DFMPsx8hsG8j8S8WkFWJfnqMDYuJiNDrgF
`protect END_PROTECTED
