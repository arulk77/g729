`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Gnmd6/n7/vowJ9GeE6YDTvGsbRdbzdd/zfAXGu1j0BAD4Ln5dNOYwFawBLF5FvrA
LiblX0hewx5XQ+t3s2xxeW6TdXwfoTrElGV+DHe41HQurw2w/NkpHjRF3YWzuhSn
cd1EtLmkIrOyDGqbevwTiGMFUYTVCfYf2IoSV+eYXOrWN5i+lFWpWMk9F3m1s/qN
2oI068FUOuoEBITdj8Vbs5BEhfviqrQTLfCln97hT2g=
`protect END_PROTECTED
