`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
qKvDQ1dYoFBIIhCySb7L7sUOcNkpLlbE15COLPLbwvF3jtb+05tLwuEA3c9syTZJ
/UPcZOBM78qGrfeFbJb4+iwi/AOVHGryAOFB83JbB5ol8LeSYKBc4s41WmoIck5M
7kD0U7SWoEwPM4ORBqWAW4sDMHCahgf+A7shItbHkUbzrN3jkB5ZhZtZGbwkRJKB
WtSR53Sx8RZhoPMlifndMQZ1rrdK4dmOpvVvMOcobzLdev13o5xg8K8R7abvevDl
NPmS1IEyjP2MOhri1X4ESTDKMCKLt0SjaKAK0Gl2M156XKO4ohFaeYQP92pXHQLI
nPY5PzVl9dIIYMvkDJ6D5ScnyNx+PnxKO9oC2Fd/hIg=
`protect END_PROTECTED
