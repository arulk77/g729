`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ6glxfxLf/D3LYrcxYabbC6VB9uRhp4DA52WL4+FpZS
0juagznvP9g2HjaYd1MNM59A5JLBeeGqaEdsWJs93YwKL40VSnCelmGeN3ZJPxo0
qHjaj9CmjpA5hVzGbyKcVzEPJ8jeIu0rY087qzj0WYAeaaMmNGK0Av13vrTO+VFL
QLxUfAyWA8xi14fhyqvBcNfnblNLGrK9tFr5+TkR3O/aEHkUMRGEgTWtM8KIieMz
EqVA7qC0GrvepvOJA9Ylcr3FBWFTe3Bvp9VYbVq8r8ut4BKbjn93rAHFOsFwYDsq
QMX4841kCxk5u7emmSjrdVVWduNL4OKK7U0v4BU5CHqVi2vkk8CwsAjspV6wVa0q
7SxwY3n4zSQrmDtgEnyn3dGPp/UwtA/EWeMjOWDB7QEB12g96ISpLms1ii44tOgb
bfw5ykEl2SgjOH+7eAX4y2en9hpaQ3pcbm/7AgYo0kyyS0qvPlYMZnb6XsUr4B78
8ZCMpmzxnv6Fbp+fmZr7GPRPWbQ2oz1fUiHdaQkzD8rpxv85PFQ4VSalDQgCkIN1
rbAPTo8DnaMVmz9IOqr9V4t34eQ+wU7cGdbvm7JR5oMh7GMmDHrAFNhDBaB+f5F+
EJ3q3lJUqTPUSxoTcAve9QUx1Gbwjb++Z2k/olBlrfr+B2fWcupnIn0DyLUSFEK/
BaZP0+ypuGcSuQ6QNqScIbCTp0aiKGEN/xkaqfHEOO1EqVk8MDQpE9yvx8+4cMZw
ACkz0uf23D0FNXgr961GgQvMCxYUCqGMS0UsyBKhaMqzvZVgXAzvhYyhs0n7oxsu
E3AwY5Eevp5bfbvVwhD2wHbQqVEqgEoBSAwMXj/rNQs=
`protect END_PROTECTED
