`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
yITGcBolANjRk++grAjvBXgctrG8zihV9q4NIan2xxH5FXZLJZU4bUFjv45CXPsb
pPX9d4HWjr4816GK6dVV9XM8FYtX+AvnEr0feXfEvqZzsssS+lP7+ig3Id2JhRVO
AI2mYT4nYQj2fUwD+75FMy/7MsiQT+6yuk1MI8YqgiCHgjl+fc10m88SXzkoJvo5
MYnpb0J+0IIMtFCSBvOqpNz0Gf5uiv+jMSaGCnue8Mcj5DyHvRRJoRebVHolQLTQ
qI/ph543PE9lBe7JI1RbY9lAtr4jY3l0NEIPKBkZqMmGV9tU9f/Mp0Z5qvP6Fq4f
JTDs6iGIA4g+ESU6nNKtz870/o5CpuOMH1PgEhN6sDo=
`protect END_PROTECTED
