`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wtHFd5mVoSUrI3Ogg3Iz8rc9nIncdufDNe/8UGe8kiI
H54yrzeCRoyzP9LponNUQ73ugw1GVoojDYK+5bJM4Q7l0Uk62nPSm0C/LiAo6NjB
B8kEU2GXK90Wh8z5X+BkOP7aVjJHFLYk1v8rLI1sy8s=
`protect END_PROTECTED
