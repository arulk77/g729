`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VN3cZiJB9f6xREOOK65F2sGj80QzVWiQWYMMxbokHRaXJDTMuMU6yJ4A5u8L5yb7
OfyKCIPKKDNh4JaPUAQicPn+z/tyhuG3kKStX+vZa6OCQowHPWf3yk6YpbamrfTp
gbQpGTU4eQVr4MQwQqa2GGrtcAO4LRz5cNf+QAjRVkb+sdyWYs155/MGQ4A5Et9t
K4vYB+/0NvlJVaIBX2V7OaLeWckPZ7rU8ORUrzJhyupaTxn1o+I1eRSeU5nly0Ln
LEeyjrvGhl/KMKrIKVftWHZaAhAGo+nBB20aD9FepUwUbxc45BwefqYqZDLt2Hqi
f5bFFAUXjf3g08nkXkuIywi53Z8e6JbiNt1IuxccDuB6Rt5aPPXos1CgDFz/cV1t
dtra2MelkSSMwtpgXCt7lQOqLuxqtgmLeo04+WOKZZbTc0D+bpVkMwVBH4lvHxg9
Bba9JDblVaZRYTX9SwnxEVSlb2SYkck49wqu09q9neicmC5Z4ms1cHF1S+66iUqo
9DFOjm+lT+p+8M03TDjlJnmrFvhYw7kf2Nde/fVQetiPaDhvdTF5gnrU/TaWmJEg
HyATIBtE0noAeh6Mwx4g6o4R0hinKNn/Mw9RoHAp0M8mS4LopC+H4/jUsgxZ+3g3
F1omCwt8v6Ja68Dg0nXsxxGpRNgPgFgrzYxA/nBtsj6mCUi5vnO2y2iLP/le2TcM
`protect END_PROTECTED
