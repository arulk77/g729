`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MsB8QtnFnAzY+FZ87+qIz56PDpnj8xsYE2CrWoX//qOYq9KI7aJdI9di7Wl9mMHK
OAaDVlx1jdHDwRumlx7ucwsaaCHZAmN21BOogvcTJl7WLWK5UMLzCSi8kpH853Fg
ZCHR0PXX8fNFP65EEYgrS1wgd6SOBPsM45kLRFEOW+WyLVSRN15Gde87UMIFQ1lr
S9+RkALCOzbCDHHd1cKSBSkFNhj4FzSNAo+XAvEcnPM=
`protect END_PROTECTED
