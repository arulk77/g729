`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFtBgYsQ4LfRjGxRXNjDEqI8yIF7prfuItm5/yF7+tm3
2FiD/2jWAJY5A69Pl/MxDSukvEB9RqSokhagRRdrrnPQ7Guxdah8elkYbe5E61ii
HExG65iug7IBqJPRGLpAzaOymMN5GiNmobfxrZWZ7/tkExmtMCWvUwNyXj6PhWxO
uGuMXfwBaTUa/wqkLM2Q2WHsQ/kQQFvazN/T/JgspNdXYK7QH+NmBXORDcoA/Ew/
UyliKGcYxkJrPd4paSz8Ds0pPKThKCWGLrdnMzxpfdYrc3m+h1iCXPcnqVEmfnlb
cnMFcW6Pm4T9AC8/cG0P82lEm1f2swSvTjzrq6If0R2mG77MyPXGVsdsRr6MxYT2
oG+P90zcATYOnaBy4S0IiLQgTJDCnsUVTycql687McGmF+DG9NNdF1l8yoU1NMVp
pX6W6GMNbbjv0bFW5L3noYynhwlXuILOXoEnnyxxWFl9lCJtlM4M+09LYlyIQhrP
OgQarLUT6083GxjehEL9tA==
`protect END_PROTECTED
