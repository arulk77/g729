`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44VfGTrjP39x/gol8tLH/dxvRHVCjKCGvP1nlIpDERiR
epmXRmblkbNzbqaR8sxv3qWSJb+98CWreFQNMInmsnDT6gVttJy8G+v/XDE7fT0e
ipcM0JWxK88Lvmz0yJlO3q19YeGy4eR5OHuhYkcysci3JDhGO7bu9rZfIEPruona
Rn7k62yJ76duRtlu63yJWuEgRe1xRkgpS2tJHCCP4vXYPPSz8BaFvzRhJqJxRoZy
0ezZVejbgqQpW/8eFxzH6wcm/82VfJQKY8aRtaVRF/WJlj0sXQ12X+xaLCupMaSd
kzgpsCGYE04OCFOx3VnVJQ==
`protect END_PROTECTED
