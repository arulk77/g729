`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF2GnEEddDj3YnCQPgzaGEM875MDCexODzew5Tk0KwoY
r22zxHtWzQ7v4cLNmk5ofNtdYaSt9YHmfK/WPSgorLxWSjgR/lu1I3uwjhsbaSSi
KeSYGm/ZIzBdK89Gf0jAnxr6NEK/Aj0R4aosG2lque3rQ8btNNm/n6MomBGjaydr
hN1n+Rmupx+G1fZvH80IOlCiiGp+O1JHeyYeM+drf7Y+kCbdbsVYN5mXrhpzKOU8
uM69mcLq7FqEOHF++gGcKRHQPhnwEPmfYELuX8vF2Sx/teVOrq1XqDfNhdvIzgDq
GT/mWoU3sMetD7Uh04Ulag==
`protect END_PROTECTED
