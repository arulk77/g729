`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C6J6wSmNm0mreRMsuCF2wBKHtuQy0ACJ8APopbzC+sLy
cyBHX9UrHr/7Ksi+jLLml5Fl2G9fDcmv/k+qf3QoA3eobRTCzltPmWKSXX5zvx19
kD3X70Zoyd+y9JtMKfjvJhT3kJDc3ghWerqlBfEeWJ95xzCqo3TKGrYlKn73jKRs
hbh84UUBvQXaVYkEUFW2D8uPF3oFbpbxatlztVM/Vu6RMIdANcXYEZ3dqitQa815
asKbnnwbCbupvfmljv3IT0NwP6XysDqWEG4pBSgNxNqvIpfVFVjq/MIaxoBDYY6/
3B4IhxY6sgxdrCmv7ZXEsQcjrw5+UGkOxa+hF9rwM3O0QwSgLdjV64nqIax+r1jQ
8jZEEw9+kLKOLjqqEP11SIESgDJvMmACPPbbnWaVysp28LgRWrLeJiPpe5cDMEBB
nLfH01CzeYY6ptX5DTuRcZT182HBRPzGwDBdF1nj1BjCpd6H+5kCkE9k/esT0z6m
4P6q3dBk8vr62RnO2BW6JLHfXb6kbrPo5IScoKdt180LXcdqeOYSRM5kolrLBhY+
i1Z9LaHMCxlcP+pAG1gg0tLe0oc4q8Z6WXxA6bnBfMKGjyEg5DDn1wZjLLsl9fhv
LAK+HCJ/CO8QCISTYUI22XDw4Hz1PHNwFf5k6irx6aqP2XsDWKA08KEMQpmQb/w4
ZuA9Fjl5zMq5nsc6/ROcWaU76G4EciUWmqJSBRoBskazB+PDtJBJofKR91EBltvR
uU5VH/kfxTjf6qLYuBkUnL5MLfBPaOdeDEGPxFCa+CQpHxjdXPjc8yrGCcItUNMt
Y3CpUe2ThT4L7d3V1IvWXq+56xHsUc+UEKQH6DMScRJVF5SBNhZiW6T19bJOZ5f6
CDJ5JQcicfgyPbBdGLA5c2uD4dgBxTI0h8Y7kHx9YpZJBqcCC2JkV/Mtwvk/IvlL
OihjyM3SB5GUQbRDWgViukVdfg4lDuZUOrXk79tV94MDXbhK5Mq9Qq4dv7pvsNbP
FBl7LkwXD84ox5PdVtqIMeaD+N5wZcaGnyuQyHtO6L6GV8JGW9jS06InqEnYV0Hl
KWpR90j7v/hmDVwhM1nt2nOw/E77QHvrYiuXYRDARSOJxQzWawcEb843bH8DQqaW
yR+j7TsaZZWbAK03gHMlKUPQpn98vsLQ4haAFKCtind1EZh/GpdbyWiq7pkLdE9c
KpC/edgcytTKnV4M8/eejB6yGXUfjbAY7qpE0KbBJBiaYV/6nyeuoTKrydaX5Lij
cybHF8g41CiyXiHwpADeRALEJ8yaxYhXdudlKNf5OxHBVZ0vly9FoVxqVlP3ZOOr
UiE8GHwzuPs/XHScPAeVCyFgw4TVEk4HvmDgNWg4WwAfhSmHw8urbdPlnrXi0Nlr
hIrDzLUmMQ6iGJ/1ogwj4zXHZ//0WYm9B5OYNZRMXdEXNz9o09gO83VHaJdE/Y07
1N6B3Ey0/qlBLrWWeXExr+q99PYFcQ6Hq9CZRpbw7hRq+mGH4/wbPga/MMlOV3IY
gp9EyhXkoJVDrIuK4XPS+uM8UBbQU44a0VW+o7zT5v8htU97rxUgZDGo4IdmSnOz
4KBqPhs64cFlx9Bi7npVQHl72a0Vf7HGpyH4/fOt1kgy3U/tYg5o48iyiexiGo4v
D3pditCpKkfbqTuk/M5TyxEuGgGEbVdK53ID1AdTKo5jbZpHbXhEqvjCLm8odlPj
vunYS860cbx3nYmSBLF8BGUZSqWz8+PT1+ZmHycBEz+gtvFI19aXUxF8X0rbKjSW
aX0hAY5kVdcce72cAEIRV+w3q6kR5noweeIGgZ13UG+DckHdhwP5teWqLfdX2Nlg
dsdM8v+CRgsXKJFN90SK6rc6JoQKiYcTzwYNLhJtxPH4WGkVqouan2jDDRobrz5t
oDhclbGtSvdV6PEKtVvv7JAzFeTEiUgxsX+qyl2/ovpbO2waXMpyL5Yjs7Ee/PFI
euphLYpSA5lf4LYzrc0C5nwoxdluFslUgcRQl7zWYDu4oJWtpTV5yuUJhXG+63HY
06Ve4ce8wqmdfmVJqqZ+y7wjYK/gPuC+YPXm4/FNxhVSdzs7oIkBxAiXVzVb4NsZ
2pS0kQwjbFYYQMF7E3YU7LG5Vc4jJq9yKR7AHDC6sZ4LQWlqquL0tqleROfFLsup
qBZeXxyrY9Z2A9vLPuVZgr9dht0luPCysISDO/8Wd+DLJu91+4Z9UrE/U43ymgiN
2LexM+IyBnRL5jbQ7zJxh8t94zV0ubMIwwCo3JYtoPdaeWTNvVRE3ww9FHrmWGF8
LnRkKhFIN/wY07sIoZN7AJ7NdKQ9mWi7TOJmdOlXrqtldCD2wjXePrL8Rc5HbdNp
jOu7SX42Yo8cR8yMCJXPt1OGFPA7JumzNMtDhhz7VTmh1cnKR8pR5rK7vUJeGt8P
dtAnI+9PIXIbdzI+So8/HKLfIGmSYihECKQLxnxY9tT14YdtKlocWsGMPOHpVnkA
g2l1PG1dkMDD3j4fduRnPB+INRUyfM9v0Fc7x3G1QC+A+lBEJz+5cnflorWirTLk
CQwTbaVzS5Wq6HU6SZH73wQKD2se6+vza51a4pig4kBBAgplhpJqtEzvjzNA9HC/
1ylCnbQhsvSnKJ7MIBQRSVQRQ6W9sbS6rUxZkSLFBC+9ziE/TwcMpUB3Xb0FD9ox
HBG1GrKoFzq0TNl85G3F4OsRHHaj+UWpcQVHb4xtTx9KqpI1DDxJVhn8XMTJKJV7
jL7ZfZgLG9aDcthF1Rrqxe29+u6ZSP9ai7VeZZrgEqii91xQeKl42F8yzr8hw9a4
Nb+BEa5ZnmcGRq6wgiH49csMpZ/i7wfGBoacnxaa11H/iVNHByvkgDNXuAikIKMB
jWOtuBIsb0UO/5gYwS4hGSkotVBF2/hfCKVs0drcswPr+ZW4cUTQqvKH+gqlyTEv
2nPe6Rtb8xnSapWBCUHlfMuUEcvCCISbDfrBJN616hFutXrw6esbeJ+7CHgK4DeW
DTAnWCfp1RqQqKj3kJ3n70vBhYTMZCEO3qqXYkuGGQxZy+HTNHBd8oY6M8sSFPlr
l+3xfWYTcx7zZePXZUI/M/CdN1j651S9hHwA4wEx0uGHmmTFsmvoq2DrFNwb7XHJ
5Nt8do4JzMbbIy3uotQlEoxpWG4t0oqyrRcJh0+pn2bfjDi6l2dyP6jNr9pyqZLp
nYPqzVtce1wBCYELGP8Fn4WPg/SpZxKe3lLpl6J8XPIWdcy0IN0UWQroikh4VJzy
bJC6rFIhntdbOLcGGmKPuIOUayP8cWjhO69t6qyJ7kX7nratn6AHueAtJ0I5Tqpn
5p8WfRY65ldMdC64+/fb0Uj4GrH9f3l2IlOKH8GZQfaOg2yFuKIv7tg2AqrUtoxu
92TVVgXJ3o0eOXAQru8aePr7ucw1QVlnTMzkbrE8JlO7/HmmLY7eUk7IRy10oDj6
ifoHMBEKN+Fb6EkksjB/CcEsZTCKr58Iay9Nb0/1woaRVFMlkLkYwJUSxOAJukLi
LBb7L6HKBDGzp+nO4rs5ZI4u7lzTgDsfCFDxn4P5sGCF0P73co5UG6nEIwYthmdH
t/Rmbd6pNiQ10Cx6SNEI+SkgtNpabT8VN+CKmjAoG7pk3CF4CFpsDDXXeHyzbbt2
8G46gUID8QKQyszYqaUTW2xsrLnlmMv0vpH0W1oAWy1a879g1Ydl3RHi6ViD3V/Z
vapgY5ns1ylAFOYvjlxVZbFaA+GxE2aWwrWwP3SC2mF72eHIbr//y6QSrn7+fTPB
xzhf9lu9cyPy8EUqVM1fPvXGqH9vp/RE096FSc+G/QnoS24hAT+yP0qps88wYg2L
LT4sv8xSqMUlWn5ztRU137w8AaB6QjXQVaQT1EckRYOFUlgQdzNcgSEWYvka+GX6
HGvOsm0aeT6f023HK3RJL9Kqk3eliPGAVsT0Y5cz+l+/JU6V/4XNWn/zOJaM8ecJ
B5KYj9TLswH4apYk523eMu129kB+P5tvRtk3JV9jLXfW1cPHz6QHjA/4GqQpvuF+
poCEtEWyFPTsDcQUgN24YU0o/cGLnY5UsTlBohCvkX0lrlRg8pddGg37EitneVkG
A+k6LpQ7qyQbMgj/f4RntTfvlaXfQf2giw3BUpm+9PhsjA4R/0kqH4KOIApTYJAG
Bl0tprnE5VUPrglmGc/8f6gc3WDfX4/MDrfP11sLRekMUhWjGNxHgpWbBqMQ8K4A
SVmU3dxCacSlIWgKFWw9p34nFX90z4R7nT++6vxvw2WEldRpqXZcGsOPStXBSCTg
ro9rCdNL+eIfSsgRQQrNIDdEYuzkjPGu2mQA7j8Q95WHhExVcZ3a36nHLJQXszsz
mrEbx8bhd5CyRdF9cKgT6oRdfo82CC10+/1lGdhfD0/D/dz2l6LLJlC5tVZvN0FJ
6vH6lVsmHvVXDJhhGFPtRJ2mjeGQ5EHTdu1L+9/3hN/HxvqRxi/yzzNudbqK6kGP
W+Fqd8lNWSH3/lDwQqzjwT6a4RBs1LIGCPvN2ccdFePxiidrLgR2OjfjRzfOAhD/
Qew+eDYTizMAP6kvOpmAcXIW7YoVzl+74LzBE00rnxLlI53FQmD6rjzB/WJTXs/i
P0d/ITFynOB2xCvSNU6TLMWGetWAEw6C08C2hdOT2gHWuXfM+VChen1mV00X/lpu
JzYqnFKIn8egmzP32mNgBfPG+i8jvOsGVX2Rjgh3YsQKcE33s8d0eGJyRmgDJ9kM
SSUpkDcGmgBwruHK9Q+QzanWyi3f+oHkQFgcfDrZeDZol3GmOmC3Uyq+xmcUykpi
HIEnj2KkWT9XWiBAvyFJ4g0jLaS+jpv7zE8F3lk+4jDL+/GE+2CqLlFNcmKQbLSO
6tLXqEqzWaYi7G2Q6V4Oz4gFEcFmErSrS1WQfO7gY5Q8nEswczdYRJ6t8bPdHgKD
NEP/mSOQBT+e02Q+2PQv5R5lQA5MQ31Gv7GnmRu0N+GTqE6NkqfRu6CeQQqknSDC
cKQb54y/IeC9RoA3/zi9k9tYJhBr1EB+B2N5Uo8JvqmhUMd0FHG10VrVnD1tEbpN
lRQuDP9QIobIaKvM2zSiPNqC0FGe+jQtPu5PvtxY1ukY/9254J04idLuQsLttDHo
zl82esVkyDKvo30VG/4cEux7XH6JAlTy0LyBVITpw99qxwh4vBrpPtUyjB+R4W32
lMDZ3d6xRwhZit5hXPrzmWinDwRZSmhYL5hJD0e1gkVbkRM0L5x6t7FBsAFuyfhE
A55mhrBBJaYcSJkPky8cZbBhvqbAjFs1ek7/wNM7NsQvDoo28zizFsx+pphNRYsw
UN5qzAff1lCdbgoqz9R/ZcHxeVRYPKt8IIJnpbhBA5KzZGHARkxvfB3yOJFhd9Ol
KY0AhTa7uvb6SbdQWuO82SVVY3mSpsG2RWTcd4bUpLm8zUFo3y+sOylQjcN5CCM3
4ixrYC0hkonLrXNeuhBYhJhtfsbbn4MTi6emkqX7knv/CI4lacDtUnSkRPQo3J8Z
N5JrgC/ve4/Pum9UFXhkdNgbi/Yj6+YYoFxg7zmpMSlmwwY5GNJg6MX40G+frOTf
grEH5wDPATYm2O3tUZhF692RzbV8trFM4aJGLxrJ/07PNX7oHviCtL4ud8mO0j64
Q4jEqxz5okBQbFDiLMEeCb4cgSpw37yka7i2I1mPW1H9fDo/ykPmFoXRafmpkTzU
tf/gDgqjIWrqoxcmY2mscJ0B2RLouCLOhLeHBoDHRnvpxZKMEMTIq5D4ua+d+Sgb
alU1IHdKONCicomeugiDFYXcTWWKjynRthlZQEmTL63P12bLFjrYKntG0b52Q0Za
/UUQGTM+sk3q/cOXN9iPvGlq/Pjp4xn/8yfXiJAJEfUQnUwLSUg+W71TOmp1HQA4
/2/310kpICHT0SgBjzm3GRQfPBFXEmmfDWcnxZpNUWOQeceAgYncKmpZCBc6Dg81
iB6gvf/0zZqQ2IT3Q7eeu10NRQu+GggEReBnp5++mSKA72YwLIdJxthdNa0WJgT1
qUX2ADPGEJ2yyP/i1HHLgapJOXWUhjXkAVu+lbgNWIDQruRL9tBXZRLjP629KKXd
TUcvBnL3/SwZ+88weaycKF3c8nE3+PPXe1KWPVw90ErvOg4UmPSrh01LvSbYwS4a
WO04DCJN6vXsPi23GdrVJuVIU2khbVgVcYjFSOo2KBO5Dz9+wZMdo8od09Wq+3uv
uaGY0UkVvsuRDfQwpxUqjv+vb3n0H7y3q/Nrr6SKcFNyVgGH/UZ36IwBQGpG8z5T
1uMXBnNOjsJXhV6gNTq+wDc/FnUGWeNzT4D0bGFqjBlq0LfnamVihUxhgyngxzPJ
UNCIy9FDHtjk1B3wAkK3I7XCyFQmRcddqINXQOH27iGvi+AkT3RCdDGJ7pQI4Zt9
ARj8ggL8lJA9jin2cySi0gzLVkpYkf7wZO1lN8Z183yuV39WisLncA3yp7z6kQzF
s8hKbXc+qVGoqk28s/e29HfNhnaZI+mgHKHwWyKhXEOIIaA4P+c1xddovEOOFbsU
nm0P8JwYJYAH+Aqb2KTPQ23H3JCPvWzjfsDpkjoxiMFsV6z32N+7YxuNk/rmx7tG
9N30Jmze1hioicyz/k+O9RojNZol9BdPX9lJlO/LeDCk9kGaKRJVbgTkC/jj8r7y
v74ErRvcTfRKEkBYCAoB2nGit/SIvRW/PezsY0ROTJLDntECBbyStsg4THSMjGTr
MxEiQkYdFmUJcObybWs8UPRwTtZDaeaP6lNmhjvC59wvRcmljbyoZARV2JtP3sxv
99ggFLmPzQg60SbccUeKVycK9sxuS40FjOzhFTpC25tzKXQfKsPtWwLMj/qK3aKz
W6y1JiKpeQ2sYtwDTZbvzDYv4zC17rr0e/GtsHW0Ig9Eq0jm9Q65UlgqBZKEeUsW
J5O7cneWFGWOmTFrvTKFA7sWq+Tjm9Ix5OTnPCul4KPmC7xSSWJOaoXRyvBHUFYi
HdX5u0u1EiUMMsvsMY75PklJqhCEQauZTfYSxZ8TWXKwkLr3Rxgryx9jjFXtqUxE
/87IipvN7wrkfiB4eslaNvIXU3Ot37UbRG7FG/XAiEm9c6pllR1yQJUwM3wG62KH
vRYiCJj2ecYhn+DwNCSjTnBDDA1JE9yMg1CfyTM5GdxHBVSUq8/jGPYn7mh4Jbec
Yvf6BgBHLFRYkTPQ2LP/9WXWb0SrpxBOUsW1uR3X6xLGCaOiLshIuiUOT1tAwLqB
JW1NX229Rv3sqF24qDhSZbnGd72wY4UzRjMALsItcslsHckcaVKzMJAs8aRxVJa8
8j/w8PaDRpz+4Jvhe0vj3eI18POWLxYTDE8ryflotLNmoMR4NARR5h46uyhK18m2
mb3bToN68rQd4VODcSaIVQCB9qheikalpwh94+GZXPr0cxot6p5N7O0rdABTCPYF
1VsZmhvgOkXhH8aHdOUbXTVDzrczDA9B43MMa8C8+qQSpYiiYaD65rCslIiPaZPl
gk+A9n4/HgQ8/Dge6aBgZ/v5bXE7DW7hPeH1z/TaPsMqh58MikDX9guYAtWY0YXe
ifmdVlQ0Q5THjhCOFG+Q1PtNJzl/dBCEqJ/FcZCCOVlGVWlDct9Oozrgm2IDlxtz
2aIqkx9kW/bRRUORS7iTS2tPkUTggMv60mMRkOxX1pNwSAsEe2KmGFShZD/DZLY6
PsBegELz5pJwTJtE3PC3rQ1Eq9oNcdNbCZ6LuglHHzJlgYCGyJP9WBehYfpLdzYN
/3FEAvJHXAHRgkbchKoSTLyJhrQ412at18PV6m5DEUJBIEfK+zKA3+BGxTbgR8dT
ZNFqL7slTUOQHJbEW4yved46HCftZVlK+nV7i3L0a1bXAZonqjHld3aLfYY9ubEM
soPlSWr0XDyFL2biYICiFPGS0aRw9YNBUx0NLOGFh4pdP2ODoUrf+8vjvUZQoRGu
Nnaw7HPkh4ziTc1dja6AF6q3++QFpTkI6Lq1ok7/Cy3vPJjUcLRDmndee+05X/cR
IYgO2Izk68V1dgNOKVgpF9XeRGhj+4pEzymJYhfnvB0SDPIV7QQUIkBGnZEqUOdt
tg88I1Cybd09M+fpOV3X09pn0N4rvWu+a7H0aSsilwX36Lq+nyAL6yk5zmQ48C5q
fF4ZOS0G/1yOT0RJbNYHpzCMlOaEqIC0PAEIv163s4VO8GUmut6fsK7F71XHJpDS
t7/qd5PxzON0dxqLqQeQinZAzuzTcZucAO9XGFmdmauufNTPP/TquJ1f3lQ36CKk
xF2QUUxCAcDViC3mR5VW8yitFxSKu/D2cJf6i6jnSQJb4IEHZ4U/QBsx9z++W72f
ZwI4edf0sjpTI49VvrOxx/f3clWtdp0EHABAmeuFDtLfh2Es7iPJYMC3PW2DF3+e
Ob3PPEE3MwxcaofmFbEVUWQWpRWW69FMuynae+55yBepM82ZvJC9rv8mjqJPWKvt
imb0RiBAvgtQPjbRbfM0iNhPl23JZuG3o0suoIKsvN0YoF5hsXIJlxG4j1J8yA3r
uw7z6d7I5NJTLZQOLE70JrOJ+v3m1eCg2u/DmHHbaCTSZZm4w9iJFi2Ut93+OF2d
LOLoehJPYvTn09h5x2MdIzV7dy21V6V+HPS8GvJBWSExQSP99GFlOjANdBrMGNPz
Tx8W3gF3oioGgwfZpJps24NH0lJxtn4GdH9j2Fw8Rv2pNUwISEhX79CWUCGSshd4
+59QhFeKhmet25/dmBod/kuB4EXUBqqzm2mg2qAYx5MoKwUtCAWKz8SPt9dMtnxh
dy/k6EDLcv3Oc7yBzQ9t7k/Op8n8VwQnfZsh3kgjbkDu/LzV95xwE+6A4vixpg6a
ePJe55SCxagdDA9WdTHzwuirNmoYGyTqJn/bq3F/QmKQkFqBHgjYflb5rnVAIRHK
QDQEmFYQz0LqNfWUG/zH6Z5H23EGBC2fMjzX71LckM05eukZELyuN80p7w1tDJ8i
XH0fCmZ98e/9q9vw+JbhOthzB5tvjZxcOt1yKsqxo+rrLZc55TsDF6gplxOwegOr
4vZXKEUl/o73DYKEAX9921ND2L7IqDjioIvC+xwb0wZN24Ymmr7myrrKuRPYeDGZ
1Hpc3oFZR1yUSAZhoMlhKw/Xj0UlYx9WScZmySv9q0psKp5+AsCzRlxV43lzjA6b
+q1nsRcNpsguHd4DdV9g/tD0O3bDowj+NYwJJ/RcyMEmBEypn3fDKs531S/fBZkY
pYvUncujnAHmy6Pq8ITZQr/xxKiaOZ2sAYONY6JazMxAOIK3vXnXmuMMQkid1KKx
Z05iL3J6MwKEXVDaZ2VMUwkpE/E9NLlsgCZPzRDB7uhiCriiCTBKe1uiCa4oCOI3
f+lPlbizRA7dFf51o8WoUpcazCnZRRdOYsRypS6WqmSEsULTzMyPZLjbw48zLGbY
mDTwfdMHZpIwD6pK9wOMeQeUtn//s+8fpEdOoYD3+ThpaDQ6p3g+YeOLW5WK/Ecn
9pkYYUF/GCJBoOpZ3E7I67tTXLTnKgmc984zrcG/J+UPKQQFP3pb8XVl+5GHq7Aa
lrw3XKB3+r55Vwib5k1Muv/7+3PrCsMCp0lFCQQslK/YrrXwX268oYAhhyzUeFCT
hh5Vvt9vL8P2HvrvnbBNNIH5NBOM5f+nRTM5l5Uhzgze8rvh9dhVgftRkyqTcNuI
4tSYC4SbLm8GixADQjBDV14X7eo7Z3MZjlM9xNLDZe0c73yMpx5f/Is7gISwBd8b
lVwwmVe5qu+TBckffMkkaCEoGkq3Vy50bhF/usQMlIBG/UpaCJfxAW2yqnvjg+yf
k/M2qZxRvogpNQ/KZMmuFAFlS4IenpQsaEaSXqZk9GvDM17bkFaF/tF9uRnc+kTv
K4KcR+y1OckjZ52J+QWPJcMOkeF2UidkCC+TGNa1RbtYgP840Iea7INUxgNwsbeD
p6eU9tGEQSv/OVvjN2jBcRLw4Ys4rDVAnTwN0xiQVlhFVgPN2dST5ATus+pGH8rr
FwT72tCYdNLAMXubRuRnj0u7R2jcNZt0kgDoALFM4kNY2zoYnF4tRapAdPVcW8h7
pDQ0uiooA+1zvwsAUftQqpr1Jm7Aw17uSHqhqg43rOOYzr1CRCUys8K1NiRll/s8
BHIplSuRq8iOj6+kQQ0xJ4LLLABc0qyLuD+jZSR33udvWsb5N6jEuBQ6BVPCFoZ6
+gn9Yorl5/d1y/74otZH9aKiWlXSrCeaqGJq56wHZ5H7BRk2+mzqk0g9wDsLFAHc
C5Khbc2Kuen5vdL1v7RqgazyRaeRR9IaDXBa9d+x444WSnfkVRlg2PAOgsM9ws1a
LtaAy5+mgaMnxiAuSEcIUTztpib+KpmlQNVfmAQX2SwLgULV00v7Hkw/KveDpjpe
Mj0ETsj1YF4HlSJnOBZXm1TIDUZE5dLmjLUe7WQJDbVKMwGEQW20gm5x0JGXSHiH
hczFO3NeqKj8+wFw1o1AWCr7eFFoKvzu6a39ZAlXmjeX1eP3GeAevN38mK414y2U
DSjaztqpxP30wOP7SSM0NsfaSuuqjfxzdTKgNTlIGDWZLOczgCCtBfRhdoQoo2NU
kApEq2eKnILFKy2GJE4YubwqNeZFqTQ5mJocAoMxsawMxqH7K64mdO13PmxWPeYJ
j/LLXFreMfttqNaPLHdbqrWSlWK3KTtuB7SjNjOaewY=
`protect END_PROTECTED
