`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NuO3fAHgZdXGyVwnz1mV3PWy1XYzGgkW0Pxna8LxvuO6O39STDDI5hz9W5o2lbR4
MOqOycynqZtUquLekfQs0SZ4at+CO1goSpeOjqOR7JMgFsbHI4JnBichD71y+p9R
mf3HgU+cLXpjESNXqdiUI5JSyFhT9XNauSHWqxAzB79ZvaVuDeD95hyjIFChl1DA
4wt/TyBtgBEWU9MaYZ6jKA+zLKhMnq+fVzguUc4XZCcXPJEqmFl4Lu3otzyQpmCe
RDaMyaC/5zWtwdRCSTO7XdVzF9bpEFFFJcHVI3c7LapznLdOvP2nbVfXBCEensDg
5QeLqfSz8qdpZlT50DqdEJ9XDw5MFaH0EPbG4WqOkJAIrH9U7rHRFgI5A+hMn5m8
6gtzMgWcsqoQ9H0rbFRhkLkzGjbD8tGxR46MJa4jZI+WLk7aTXmDhMNA+8IDQMeV
1hy1Ll5A5Fx7jyPByCNCo1noQflYBuUEGrrrAoxP/xrOpkhEQhbrDsRCPT7UPvjc
Y/YLgfzsqmc2fgzmCyMEi37+pUPSa2FzZIrMPSFlltwFN8kxGaCxMC0QDX1jcJZR
dwT3Nd5Cl1okJiYTyXnErA==
`protect END_PROTECTED
