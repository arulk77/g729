`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOKZBHJ5ttrmubiVTnoMXJ3eq4I1VKv6z1oiADa929mD
PETMhU0mKOihUQeHzILC7As/xdwPjlPXhuEFwzLILkmrU+csH0G2SMzXXgXZNVW3
Hdl7D4XYvYsIxEV9R2vfMTq48/ogWRBN/tV9sboLAg76GwdBu1Nr17QyhkCjcoZu
L5G8OfVQ5IR8na918B7tMPfOojRZuxT3ju0QgLiSMnIxbaKM/irW10PVUnY/rAT4
`protect END_PROTECTED
