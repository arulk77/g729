`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKFr0Zliz//YfR/SSviL4Hq8SHUkWdsKx7twdcnFNP9W
PVQ13B8rvM/O8V9FVH6GPiJY66sgEbF+KSz10lg7BToHMejShzOri1Lt+pUJNeNw
UiiF09HuBi3w2FzlJnx3x/ERNLrFibIOFDza7vhWpQ0iNs/Jrj65Ug0d0Q3XznUc
vl66en/4JzRalefNsOhkUwn4a4x/zM16+fJXEIOeX0mOZuKpUa/XUAUbJpU466Fl
JcyPq52MSbhjV6fVic8oVgFyehOp7r18sRVUnkcz3QknBfIAs9WuclBs803pXZ5G
oKCjKrLTxeKpEZhP0QSlwovJtr5PnxqdxIE41vSsi6eunfP9iuv7SdhJnAzuGzB6
rAYVtix9F5QS20imPoN/iwrVSxZJSYY8xmuKz3CN77q7rvFsY9rb5mQcYwp/ThNf
SyCBEUZSzirEGH2/vImpierOrOBaAiSYC+REARde+F+UqAtQU7jzhyDc/WbfzHC/
`protect END_PROTECTED
