`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAUOAKAHdI0HrR3TdC3VinDuF5Qx/PWMswXA0dj1EB0U
YG4/EKSbjmMnK0BK14eLggSrpiUkQr1JAuhivNiDofsl87+lnaggUfCdA6BgMkkV
gX6cTaTCuPsE5qYysE269+mim4Qz2AsCkHkP3G9/t1L+5yPLRGyofblAK9c+hBzi
kPZQwmIs1E9tZJAkw3OzomAImnKcDAdkkoADZc0LgeyfPozrZC7UNa7I6TSIWEVG
yaPf9SobEU/r9qTkTkW3kdsWyQwWOHXKpOIhQ4FjAlp2cBDGgpBLDqcRJlzVfNiP
cT1E1oIVxnXgbZvG3zwqkwCtc8kvAyWLrHHXt6mWetWJtmXRmMsrdYC28oT66oLS
Nai0AakqWCKLkf8+vPyHow==
`protect END_PROTECTED
