`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z6cdZWelNASwefaQLlznBtatZQ00NgwrYq+yCCPdvfX
/yKXfgfB6JhQDo7XdO7b1+xiV6hYgoeXx0R8Lspslq1wA9Z4oGGFKac0aQi0WdfS
8IWeiFh9l1khHO1cheqJCdBmcgEZYWVYb3+M9ycKz6ik8f/WPSl46VU27QpgHLUO
k8kk0vWlRkgX/jJz81VE7dBMarHeHhUkBmd2BaWmn4iGKq0QRI4/MbDqVoPaVdm+
con2b9Eg66baKCbb/JYBBg58ob+2c29UWwQeJSsc5HNV9H0p/1s24cCw7ooL3aDi
+G2+MnQbTK0VkkSvRI7bFg==
`protect END_PROTECTED
