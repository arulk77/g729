`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0V6Cw0gdmq3VqOYojEpo+CTlfpeh2E0HwEKlqyO+0sU
csFYmHypaqZIrpilqGo4XO704l3EOh3PEmI+ZS/41JqQIpa3IrzrdsnSRPvaVpz9
15ev2MEDO33Gqbjki3S/1vVL0N1T/8n7A4/UGK3i4YCWOXpetP/d87W8f43xOJkI
4I9KEAwd6vcIo7jMgt5ADhLJ6FonyBaM3S77muCj7IPVXyt/bVoV7GAk8rS1c1C+
WL6PbEsd86in7oOZQmZSokUCeaeXNDoBswqtHx2Rn3IR319vleaCCKiBNfEtqM3J
m/LElYp0yYJgKoJ5lXEmBv/ED59Ypm5Xbz4uIKDwDtrPDPBPegyp2dvVJbS2zmI7
sIXsctXL9yZrATJ1zgz6QY+RDKdBSAyBBlUYSnvHMIp4HnluS+uUDbsqQU4ziNP7
3dgeOarUUxYLRT5cjUXtVVst5NFQdgUkONDCTrirKc/d98NXTzqacT2if+y4ZNqv
LOZVTmMRo3w6eq6Avl5QMcnhRRRtOmXQsQIu7nXKa9J4lTBWClEaISAsUWYuSuJJ
NQXdU4WRAb3Zgw8bQLTNLennCI7uh5ntvm2ZEIEG/Fs273dfyezcGP1ntv8sHo95
gKFXeRWnfGoSgka3o/mpi2+DkUBhQOmzQVuwSFUrf8gHPSEtRPKWqk2udL3qbzOc
btbfLPKb95bvLcfWEyRRK9gCVwGSBSINYMCX2GYVedv9r+KFcsbZqt+6TX/tKgSq
xOW6sePBXOS1wR9nZTgVALZ6BsnW339B2Cm/Q17eitmNkGfyYnb54lvlRTf5zACD
XvMx928SCYJv9Mx1uGTYZLx+DtrPg1bGde0hRdjD8Nu+mYBPoINoM2KTHyNy35Qm
HJoxfAi1dH0kqWXG/4L5GlBQIQDT8J6/nby/KJdESgeUlPw+L5b1FJMv5DxK9Fnc
YVa0b3ufp0+uJK/M4+2HeIMJR2lFWWOlrdjlCKQ+MfhlvXZaZcag9etU3Wh/nGcY
DBr+vS2XysmNjNKPVvdo70vKmMn9suRW+6Lgg2Eu1phGWr9AtOdONWkMDuk0F7ze
4PHLoMm09c/KmTVsEGefZjNGrxs5T0PC9X0vACAj86JcG3jxsbWN9nPUJTkIc4gG
QlnqY5s+q+sW7nlBogHeb8KYKrX1pogmOw81q8RYdep78P7NNUAk0IbnAlv1mlNY
E9oo2NJ0NZ0W89FQoAx7dGSl8oU0LDKaLxy+MuZ68npccax5YKW1pXKs8mX9t7j6
GNuhCpRo2jfus47vxZx+swyDp2A1ZBj6uNxs23LWo8FcuRogPtIxgTXFjpK1e1yx
qpFuBIwhqaCT3krzUoUZBtKeLZNy99pgyP/qXFztRLCHN+J9RFBIhFMsX4DgGpUb
od6gD9VVFyeD2v48IhLCIXVc+6NRVneE6goYsfegRgFlRVpQXwIDDcCA5xrE66R3
MxsSqTdgEpKWiZSFM3d6d+RT6XX9rUKrnwt5AB6vxAecnDN7WX0M5BzOjxXZhtmd
uOOc3bmOFgnxDmVMa5XIGI5TC3oWNyDbJvnYd8NOrag5fncEzCnLl5myEciw67D1
fY3QT6qhchbr3tpIiauN/ZEamU+xgY1SofllruEsvpi/Q1b5Bc1MWz2UXvjScf3Q
gOQHwKnf7tzXmUrOAwpehr4qQPsIzaVtWdf9gjLErLudVIdQzIL7V+PNtNq1DHxy
EM/MgypMR/M0PMmWyoYPdoaqLDwDC+ROHUSEbN2yMS3g+kF8YXFJlqhTkargI1B7
/DdL+Ivg+aMyOFT+wXUnQpMEXLsnqMqv9gCbOSmgVLkJfIxHgyESaWijkv1d/ldw
AYc/n2p5Ya7okJVfSwozR/1qfPtUdvGJ5fEp3ew73yTjJoOnLWrzxoUSoyYgPLMV
aslFueKLHCWx+5voT2cFDpWJHsHtfO5gFyUwQBx3absNxfqF4Bk+hMz6kky2DJ+g
AYBDuvgQ2Cte4pWzRz0Bj6iboMrPYsNUO8V9p/TWduOCpbVGdNSDaGYBUHj9WPv+
/jWWdmJOKOnDFYGWa9Mnm55bJP2V1sEe+CTQMHX3dK4cf5n7UMhil4KfTaqIaPDQ
RStuq55pnshEeOX0pRNp4lClFvalNLoYeUPDIb/EnWYPI1oX5ERmnlTd7PM8VxNN
mX/1+5yDXi8wkD6IDDaQ4qWB2aiFO/lAUL0ZR1tZrE7Fu1EgQujLD5ASnt5Po2aS
USdZHb2u+LWgGg+xdZPSM3HOpk//mninrRMw9AeBIiRxPXDOjlTLI25Smgv0YxgM
6NgF64UvnW65AnwuiFqo4JSR/17+pKo8mqHc/i6FQ3R5RXboIZAayIOP6H0JKpVa
K1A5kM3U20Wg+0gcJVMQnKMoyFACPXgpDpEwIGLzn2bvvoQEisu+trvxDfFVkfox
MHpoG235ZtaQcrShFBuX5A8DfktQaFOgRli5JUXFvfzo0PIPBp48lZO9s1s1VIHJ
RHalVHPaY2USpCYL094n9CDE2pIkFir9o8PVAvB+ZJo=
`protect END_PROTECTED
