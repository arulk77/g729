`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TrCVeMNu1qm3rL/3Ol+kuEGq8+NPROSbynuCXkjz5WePjDw/AVCXA69IuKGi8Ov9
D7vi65CI2l7kCUouISaOpA/CaIilRaZuPOk310B+KJatlrGuCM+12Rg0vw6N0C7F
GyAS82tN8k5YSA+M01qdVh5jBjtUhGNNMWAeLSKfrbNF/pPjmuCrcvAL0YiVEDhp
m00gzcknNAo3DIOJIPtLsRcXk/PfkgReqWi68lHNjNcr0fCF02roh7C1OpcJw5J/
dakUhuK0cjdZfYocqFDMAjoTWbsz+F7vRqyDPfoPoOs1htIHGhbwhMZwaVPgEBPF
d86JjTmAtL6ybZ7vZalG/xvTi2YhWI4/YzJFeArHDHw=
`protect END_PROTECTED
