`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD0YTYZDx3zxG9rghHP86on3B62LBoZL7C9rg49LezdI
y3+2+6XhQfQu/km5Aown+CzFzHMq7RG8bIGLw+mJJCTq291ltFrERMxfhs0J5Dci
588+JQULXJzzyELguEHodcdkI6GKswgurJG+TM4Nn9ie5Kpif0ZZAsvze3Kzmr4N
DkzzjtlL3sgCoqYsdOsvln0vmAXegkwqM8fKAGOU76P/tTkQR6bwcNIb41pbv6yp
cbwkk+fL2C8aI+gna+W33cfY+gDgE5DL2XhnCgYDCUkaLW8JVXfgJ8tgNhznL+NH
svJf8Vhqt5ScIRqP/M5EHw==
`protect END_PROTECTED
