`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4viP8MmpUZx8f8Mwz0g8xdvW0lBrnG56TU8b5OPmjBsAEXaZCEmoqkqSleJw3NSm
RsgZrSqrJCNkl3tgut9/wnH/5qD+6fqMyHuNFF3WjZ92ToPuGagst3eiWxcnx126
k8DEFaVCznhWWiV1oL/8yl8tZ5WLxuNYPgpCWksc225kV6z5ibT6DXkfYrLzLKCD
yaR5IqhHFsTVuwgnYFzTJkU55Q3vuZAt5d/M3g8nSR7jAzjoz1Lu9VOYZzhuLHEI
gRwrQmUvzN+AvgmsWMMf3g0Gq0bKKfWMFr/nBMM/JZz+GzccbXj0nKHNzqKDWzQy
w28G8JCNk0qkOZZfYFgvm2JrD/I/0Dt/fngsr14riHdDvc5tZ39YGcI2b1+nEJUf
MscPQ0rMdSMVnKKtHV3OrDjsJ0dwQO3PP/ozuk+EwZonj0SLqzm9/1GDrr9X+hLP
KBnIg/uR4ahwADqoTN2I+g7DoaTZYZAdBtoMNeeQzGuw70syjYNeCude2T+kDEJF
z69dyfMq3qmnUSabjPAoJot6vEHR4PtQZAKUXni8TMC7G49tYA9Y4UZ0lWe9sIVW
4gJVRoMY/R0CHDYx3X/kNKZB+kGoA7Z4Z8mdr7IzjVBMC4LtGczZimWuz9rWbkiT
hvFDT+wLEXdoMpRhUtzFLh8UR5TRsEWd2LRQwcvZhGzc/phzU8sZgmun3P80dxCI
U85Q1Oh0L9t1J3wYEO1Eh1iNlkPtv+qwlvJpgtfwUUdXT/N2P6QXX4XC0RgwB2B0
yvrPWIwgV6bp53hergrmN7sh/ilML1WBxRL8uIO4B2gXPGcZQVYyJ8U7N/bItyS2
QoVZrt5gsSHTbGsAMLFkhPxrE0m39Z3JmpK+tzaEtEFnyVW0w1a+hYqW7/+3VAep
vldBsCk9wwchBVfHic/Tkvxwp337dP8gKApOKGt9rwCiaNrY0gDviusnnrL8OYLa
bnznX3NpzA8sInvTY1dJc4PRuGF63NhtlXrZ10B1QtavN2C3U//9cTkXijNhEPel
P2mT1DfpaRLtdem28WEP7T2m9Izzx0FiKlraHUkbEXywRrQZxQc8hDajBTTvShZ2
vXO2Nd1PB9iT8GwiicszNA1yn8Uvi6Biq3u3BU3+vNwyP7d1r7JGT7vzZGmMSvPT
VZmoZPaoZQuxrL06dJ3x735sDYlC0VhEVK+8CKHnAhspIFBJ3x5Z7E/ZeSlLlkUg
e+mPFjoK6f2fuRgbormezLCHFSiZG0WOWY8f25V7Hs8mVWJgwy/3o7aG0xLOcYX+
wBzNiXxwEc65NwQH0IKpl1MoVLeNm4twCTowVPvqXUURiXEoLSq9EJwFW432WYfS
Xnj95tfPsbyAaEPdeGpXnur/LzGXExKvvWjxiUix0N/2ZTWFpV9znlJ0qCsEaytm
J7Dv1AOZb6zcAA/3S8ag8QJdJ1Mkb/nQQSpxX5oklL3cm1z0mgusY2h8xrHEZUls
nKesenr3DpvWlEXwmXvQNBi/rufYbs7smN2jVEWy8Vu5LLXooBJYWu7N0l9i6MEy
kxVHOf0YOQse9WPcWtn9hQ8SVeSiZT0d32N/5d1FOPqrub1M56WW5YoWwDGs0XQT
noz/5ARnAry3d2pOPynltO7kpzbAPt+dc+wT34tv0YLFjhDWjVVAY+ZiutT0hzPV
7jNHvKGVMix33MvsJJ1dMVMim22GjGabYJKiZuHxsXO1ZqG6BuVabCBwpvDs1pEr
qq7AmrSMKFfOBHzk67MsJ7xjlfrs+9o0ake9eCug+GxhIbF3tksHd0J2WLXm3H8N
9GrPc0FRYPkHwIXUKeQ6WNFBYdo0sYBmMv0GY7dAEiJe5Nh3//r4jqFZ6mAgBcO1
p3zRJvKkOLdG5kEJ4kJWTgygPRO0b0CIRGso9oT7v0RZRQsFEru7RDrj4gv3heem
Grf9ygn1bmLM3wxC9ErWZL1D6RvP35zPMgHyJX3N7nF9rl+A1Rj/C+fjp2p72sOZ
EJXd6VZ8tTPvK0VEoVgf1xIujXdLCNtxdgjcQhlGCGdqT99SxaIxXV9TDNvlqufm
+E8/hzNJbL1rJc/ql5ngXSpBOMVNuxp+Pimffkg5/M1RHFmNETpRCwZ0g5CjDRW3
ZY2WW4+h5ybMxusHdZsxokX2hNQulirmIlJnQoPM3i+KpJsvh26P/R3xJe8gucra
JGuUGB6B8VIPFCe4tQcpoJCzPjTZ2ySvGkTkpkeq4o/3XCEnRzXF4vkfstbYFqoX
FlssARrZC12ANZi0Ndl2D9U4YFV7WtslOq2CJcTt+MGtbho5unfjDXwC9ltGFp8z
THWoRxk7q+D9KV8Gp0tdFMNK+hlrhmJ9v4kniu4ZMl4bUkCk+D4wmj7GR3oLwIeU
4CNNwrGYXWIV6ssmnOi0kjGKdv2QVsOEzRpv0NksvHhVyx9saqbdME77gB/YhC5U
O0mToCp+YBvQzZD4//TaW+zTaYSIeq2GUiX0moRrllfFYBek5lGlEz6J85R2VJjs
EacFfY9dq8e4YFFV6HqUgDWS6UYk/IoeCuzoCwziZo4dg3DRwvLCimNuobpieXuN
YWo/SMX2eY1OkKwxnsLsvqO2XFSWD//BpTn3+hlh/vC/wuqA8Oc8eQNcoyzN9eg8
x7g5MMq23rfJLG1xdd3I0QkFDF5Jkd2e8SYN11tXtUKJuUuopBpjH8XwdNTErCB/
B+wbsCCbDlFU6yP7eCifU+xtxvViVjAQZPXcx3/0uUEeQSVMc6V73iFpX/JHnoMw
1K2fbp31AT0aENwMc9CF2FtN+xEYVbCHAU62iyLOpfLf1qSRkamjwbqi8NVIzcS7
DfPb6LZCPGi904TNnq5CzhibDDcJj85F2l1LqSkC/wYhqqAFACvKMQA2q/K7mUxT
NJG4KRAvgFOU2+Jem+d0Ktlt796OrW0HyhvayAKfBO7XPrgBk9z1xp5nCetE1ITW
BGYjKA5qjl0GhK50pIEaj+KytsTxcphCf6qYSBizpkwUKVVlB3OB5XgZws/1kDBa
5EF2qNpW1N6AUzTxFp7RL6xR7M1AKor4e+1BsQc7uZ/8761RwmyhXS/hhZPzBQiQ
Pv+7jJPhIruJms4ahejCI1UNgeoVJKjRqFPRUyiq06V7EbpGm14CMHIbv+FuxgpN
3csqPQ1g+5pFuHyfuZ+nCRQ9sz5761MfgMQmUOSXZFBtePjMSk6dUApp8XM4/Y4a
Lk+vXEMEhskc5JK4J/lOGXj7h4BykZePVd7s2djVKcbdya4x9nP3aLCzaxitcVS/
AY3oeMtrsGHd5ttcEWEh+UphWAwN7EPz+nFVoJo/9wLgKfDwdoVN8p2vBeSMXH94
77dXddE1Pe9nqkjIqL65tHtKK9wCxwGNmXxFD5+fK/pJcY2UVDpL+oSngl4U1PTT
DivLnS7Uif+RDR0LSDRYOVzHHS/vBifhrtxXGpnjRoTlkxVCbQhQwl2fyST0uWwk
dD4TEC58OIi3MQ6/JEPWtKPJSApODQa2Mj2J0/AV4pTWtjP4bhA1Od4KmYKxUhPt
POgXsSL3a/W88FOlKOF99VF6KRHnKnR6VPXcmLJyM+DAaGl42GJkvxoywMI85ZjT
lU5QNXXVRJkkbtdwz5lm/k3jUV05R+VC6pQehWrzQZ6cGB8bRKqzUJVAlky3Fpw1
MPFDQmh43Ad36DykuBiyKZHOumGsTVGvUKvM+b+c6O+nwqcPhP0TUSUsVuREvEJS
z7Pn4tc9tB5dkGPGl1dBZav+4jyREbrE46m7+zHMImemyYR5b9DKKn83/vNhs/Db
27qMLlqvPGlWwE1uZHAWYkZccVku6ViFGPbV0aZpCod4WUD9PuiFY9lUEhJHtZ6S
1OiYNRWR0CZriXIPU+rBSesSmTdu3LawKDXaBwEzTpbOADzeTmwdmJY0xl/Frwzx
unW+6ACwKvtqazTq3Lc4wLWwWjfAS9EKdTFuVchpJI4HDZq9B8eiTEpak9/TdOKJ
7UQL3zqkS/0KxIpCE6wgFQqwg6KBXCP7uePk+b4v+qgs/gQJs3y8CxCGIkmuGWk1
0LCPLJsF6/qBuMtONmy9o6oSQB9vSG5jDmioMiA1EkhZWcDm7ls+Oj9KU8FV6fgT
vQrqvkzZq0+q1oKUDwzAJpIZZ26VCEYGKWYBtto65UAe4EVRUpi7wKpCJlDY22bm
LonW7vYE0OrVU7K8fbXNWwXwCSQUZ2dhw7+uRlUg7a2RxMzoG/qAQm/3Te2YVdA7
50JslB5QEkESpTJhSuuBkfL+inXoM1AX6SEOyaCnG9niykjBnghQ2C0kYc6fr1OW
sCEfOERSlN/GUpUV50QYrH5st+W7WUzcbIlhhMWynOxQ/XTBLog/HVR3UubFexDf
rKDf9nuNidrp0J1/P/V7HmyF4/wSrh+fKFQrCcbtWWt+U8caHHwrGsJo0BgidR2H
KCLGXSCeLsE3Emtd/JJOB10XegcLqoQn0M1vs3VlaT7KegSN8aXmNm09Ga3HGgqD
DQ9JgKYhy/TJA7JdPXZA1yZMtDF5G6LsDf8mRjMar37tysnIXrX7hiJQowJHpHyt
GaWuStsPwR+AYl8XESoB7aMddltJTqqiQHiICffOLcAzxmOFhiqh+kjUgIfHjZAL
SL7GKcpWWbqpkUe59+aDGc7+aJJLXXyNxwAOFegh03A0m06whSF1SYRRrEOalLk2
ZvOSL10t68lH4vSCsKurKGXHdD+I97ePpGYtA3ABaxgRPmlpphSmiTsF91Hypgca
kM/ch+JrG92REX2FH9H++0AWhrl/x0pH5tHdO/QvQQ60147cu33Bh3eoStE3/nnD
7mdhiKrtXyrjzPGJF7/FKt389ogK54ltEKFr99XatfolLhUyA6xGamVwZ9ybO3wC
qRyEIQYdgV8RtxKCR2in1/FXn8t6ALRpQrVtlFYjmfiiokFdR4F26LLz2r7m5e3e
tS+8G3/qWCaBh8eXnnsOe2gscb/DOTtW/4jpZk7VAVOL/Ii3l2gEUCWpOlPp+Qz7
DsUfP36UVqYBd0qx83dXUtpvrWiIosCr2LDW/tQ3DcqzYd+33z8nnF+2VIZveTTk
f2nAzA/TP4KEuzr9JwhXii//u9bXt8L7FDi0yx7u12DWCjNvxwV0amBeZSImjAmR
+s4Wolor4FCqTei+tSaleuiOcJhBNajUDxBaIwSVSm55ea1eodpQz7NPjwmp8F9V
5lpfjeW/5B4pcrUF7CNU8Ug6pt3dkQp24T8GXp6NrMb+3O75qp4kw9iJyfO4pzw+
M02GY43uL810lRmtc2CQ/CqvbvNO+3e64GDmr8mX+IfGvO3XsTr3xvmuLYUl15BM
59keVG2gUdimwB1/jKN7ahi8VvcH6F+5wK/8TUG0ZS6daAmtEldHae0ol7TJPXun
cYrrCiFRXht8Mbvz2kz/0Q2DHj7yWXou4QKRUHHjrJaPFxhQeRGxC5UhsUy7Uwj2
rgixNgC7Mbuhe9Cl/Q4ybKo+3WeO5TP0M1Yxqz7SzK/PR6wihuL+po06p3kCUmWj
JuPCVbyWIKd3us3/Cjc0QgLBzgqbXoaxwDBhYPnwt3OC4GxDftecucGnKocQL1PC
PsPymJwNVkDiXA47b6Rn2ML4NqqVtqCN1Id0FfcK6/r1zS0GH3TFTvvDg+XsxmBo
mlRgCjb3XezKAPf9zLW61n8RyZBD1B+IqDoxga4CDt7Kohe88HEJYSHfWIRKo97B
29XlYY9iC5iPtidxaf5mita3cDL7VKTKmFY7l1Dxc37OL9S+3zl5D4rCOlegCqY+
2PJSb39nG1BhiZDLw75eZTZ7SiRnUKoJ6Nuu+6O54z3oTh/Y19ltmKvBHS0NpxDM
/HJFludoNoKySpCbrIxJQocYDCq1D3hUM8nJGSeNlUtYZUxhRhM4IPpf139mklg/
WgruChVgpLt63Xt70UKomvu+m/WNUwOubGQ67KjV1Lgy7Hv5f9wdcMjwbMl6gNOc
wIkNMhOrUNVrY5OmvAMjYrVDmzfpVpCVFqzv41Y6/bhrVjJU3VBj0P0M2Rf+V8EG
dH5iutjo0Xdte5rSBGvsLe4D/S4Abza70IgKnGLa80TaRhI/rMCuVPd05xd1qBmu
HO7l5YmocAZ9kebRnG53z3p1bLuAV/Or9fW71Wj/C7b8oOiNKowdwsSVm82NRqVH
/YkJSj9Vbo0wm3xtKxdaadYNdfnSh0wT+XXJZdnhxX33WfXYSGPXtwyLlF49d21b
SiO8gXaLs6GxqnQLnTP9/VPk7hskVMN427mHh2+pd3s3tSkn9W0y+Xi+AEazyA/j
dvudebtOXdm0gij4+l+PSj6Ff7yIYo+ya7z+u6bhGQm+VsqRWxpAtzWfAzpKxr0b
FLLmz/My7b56yzLr6C7gQcbo29cUzmK8qX1bgap/ogmwLS6VfOxt6rB10aFQr5YP
HxpH5mvUXJ++ef9ZIflKHFFCyKVHf4I0/n8OKlOa1+v6o04GNEXibWzsqDOr/Gkc
XS+G3ZmqDI71kp72DzaQpeEP3l7LaraWhCTrzpGTeAZORKl6FtqaUbBMEZ4o3gsu
Mc7+D3yW5EfdjF65CO77tylgsRxiTGZc/jgG/k10lf2NzoOq3MmKbEluHxT/hoqT
w8fySVsidiGv3oPfSDNDcqf35bQ9qX5HpzEqdUaNhYdvq2hz1E32OW4ZlZCcjDhB
lSgvoAfmYLjICxbYUKWYGXHOE+ylp85aU9dtYRWgKfDOSO/qayLFg0y9eZ3mDodw
/xB2Usbt+V0QZJABrossL7GRxVzsV3K3BrF34033EULS1wcjJytXcAJThgYRXchh
lGd0WQGKM3lf6HaaGLUBECaT2GcWt0msk/G5r4i9jH+JO3JH2q0sPzLbnvFZlD2p
v57sMUv1lefxqNqAZnIrbxPZVzEPBGODd8wnnaCCDADV1EJVaE1vDlawkZvGy9GT
JrELIHHfT8GSVoYE/slLeTtbX5p9ZJ+OH6PwRrytkRWElOQKs8QmhSsZQY2bkn0N
DyOMgKFkbC4f+D1u5mfmCjx+pbZfM9611rsJy8V7SaCdQyy7/7bymAIz2SMT/oR+
rySTtZeGMCeYD4urBHsTyRvtX6St4E7rG407Jdq5iTb5DqPP9m/HnpRvfGKm4C/C
GdLnV/IMVOFxySioVzD4xDHwjLCswgG9GYALr3PEiJ6wuhFi/dqRWjnlU76WK+IE
YrEQacT8vaOiutNbeVGZtkRHgUc2qUk/Sa+WBU+SLnHWE3TbBdiCs9lwRY91SYJG
17WWmbBJU0iv9FVlBo0aOQ587MEcjL/ybCZTnWm4p5J7mU35ksB8Vt+n6za9zU/o
dEXxW1uRhMj5BWmrnn21GZ92zaP82Uxot/8En/awM/NwC6ZKpVBzCDoL6djHmPJH
1YwUPit+dxHyrGZwAgycxoxRKueZYl+kbxemJnrQ0zCHNQPyAsTKjgIGWylxTkHi
YCJ4qOjIk2DXVcuBKiUOqL4zBeOnqahj5p7kcpA1YvosXyOd2k/K2TaZRLC4i5kT
UQxfzwBo8LmXGfM6Z9HfwhX+OJuTHtkApzNL/Wl6rsO9K/es+Ke/vPo/6NumIrHT
u9axw98G6tVayxFVRNFqusJyVgJKhsYB0VoYUd0u1AGluxqVG7oF8mWE1PQd91LN
RIWr1le+XaKo74Ko0W8SHCaw1vb6NL3k1UaFLu0S8ix3Ka9fU9ND12oRN01b5bE0
2npWEL751ABwEGxK7jf91kMB7Ly/HYuz3gKshtITuEFYZGlXK+ALa3+OsNuMdKz6
F9lFpv0Wz3vuZXFRVDMoxDHfL0Z2yUvXxrXbzw5xa8WnxDQ2a7L1wNKxKSCR9qUS
s+Lp/46ehLEee01HXUvtnEPzF5MeddZYeQ/XF6pMuKM7MdICnvEfJnxhdSXpWnm8
a5g4sGQGY1HIvfg9a5n/8Bca5suk2q4EvdsOyq6Ee+Tzk8mb2ioBxA5f32Vqs4d6
XcbFHIbRy8y4V3J4h4LyGEaQ3dYXWokUys286qegShVdbMSjLLUz62/x3in75ot6
R+Wx93ngAMy5NN5L7Oufmzy+SfyJ2vGNqD6rR9ppY214nVuT3z1wjDoono8ALcZv
d2h+Tv2c2eIdi2G/ZYrNE83EuMeje0NzdtajgA6mg5VXDSqVQCzLwkgtTB12bPNx
S5EyUbky1ImOUNWmD5bza/A9zpSko8wMJLITam5opmtnma4VB3iMTV6BVLJw1XVJ
vs/8TyCdDhip2lalFm/VLg/mWCrEv2FkRk+0i2UHwj/jNGdu0EtDvRB75AEKQC6a
Fv0u1kVQ6LxXrDB4NNAjbBn6DHdpRdxpDAqvNO6wF9QUYoQvq4esjiBSR2qgpyuo
oITPGE3v5KFOw3TYCpLRpPs1TzQUP7wJ26QxIG1LkF59hPQEkGfpkng8kV2Kt74v
x0itnCgqQtFZ2xNZEgxZ88ynS/RgmmWqRjvzKvZkNi+z6jhEOUJeO03WhK1S3Ofx
gOfAK+HDvtenpgB3GIzanUEEJPp8656qSCRrWAyOI6Xi3UB637tBb40PYbhUuhR+
IErNuy6aL/OIP2z1M9TDu+qhtWO1YCYQMQeLQIS5SsX+2vcQOdAwJBh8f4OBRze1
OvFQrlcWQqE18x4xhNcS2O1kWiyoMa6Ihpe0HlX4+fHv0mryOYj8JBPQFQfRSS7T
OK5CDvsqW6OBx+r9BeUq8vm5UWwf5dI/A8ztZosOeR5Ae4ok0HWFrsMIkVEGuh+x
lnBavz5PpHQQ13Xc+5aiPAH/+tjkZ+4F4jO8a2clEyab6ieP1qIDje0E2aUVn3to
cQPBAUYr3kIBPDEbdfwyiKDewLQpXFNP0kn+h+0AY4qwPENGfaMZ7EA1awcpD4uF
5ouF5pUjgF1bgBS6w9d4QextTfG5wr31Jou2I9Lq/e9F3OWW4pDQK1Ef0rwtD6G8
P5kTd+VyDkekdVBrF/sgFJoqk65pCfIeVxJdK5DkQuLjNNmsd9DuXYGyP3z7npEc
V4mXmemj3ILW6WV3t+rZzezxvvn8V4oyhNvZ0wopjpFOsmoSyUKtELJHv2v1Ed7Y
pRkbYy26v7CZudRZpr4CUTtgduGHfTGu2g14YhPXWbtJ6y8ifwoN4Fueejtwf4j9
3yCKlYgXwXw7MPBAz1WQehO/e51crNJ6eK36fo9e2OnrASKTTIcI8mclZ8frMrC5
bkGB+pwXbJbOB6sru3EEtSmC06ss3PjmnfxsAux/C2fdIL1qkSiNhwu6R4Z/62V6
blylmSG6Ceyi6Ucz1gBglslqrnUQ8chrKr5iBHCHEWYBgYr7+D5TXL47pNbTl+gV
gqhLG30gfY1JlAAt91AqBplZlhsGTIPtZFEhi+AnePD5PnsYOWyYqKiU9PYplxtz
Y/jmgRRcp+6QerFDv8loAGGnNq+WkUeWBKYz0gH8jyGvrs3nu4Exu+fjmyqsQQN9
rdwxEJdn1VaMrqo6i0epjY8SWDtIA+7a4FqAf6vz+vcph0ppXOco/xYlITmUwFth
q/wzpMf9t3ykYujrHE1+aK6lkvT28UYjOVry+UDpQelLmOpkFEXMmctFd8AetSm4
xS1/gfhUddXhDdt9k7M5DB0o0qgO2uIM0Anxc1W0uhoZmXsmtrKo2LFhYNoxQib5
AoRXmVeOEoFGCY3yHDJtHAJh8B7ryztdR3oZ654thYFg9NhEgqmF6yVY55qYQuy6
3ZiVH8qJT1n2GWmhHuR6E2conj5WkodOgNuuXmjA9WTWCzE24qyDx+XpufVqparx
fCazRwuTKwnCqGAqhllnHOwrtAbF456L/cS43cZu1JtTy1p8THqxhXqYm+TooUOv
hgxlkm3dwSBwGojvX7G8BBE1GNlK8l/BK/GrjP/CcJ6uDV3uepFIDnEN0HVbQk5V
xBw4m/+bqezd8cEb/muvrwwt0FTA/f4LPHo8VR8QktoQZ1v7VTL1WF931auAoP3o
/K4zJpLOP27Bb8VTUkC5Wa4GxMQBzuLNCR1lgo21o97MWo7kMN+5ksattvFs/4/W
1V8+GroBqMv1Nzw3sQG3ZP6i6DtGSnpePwfspn5wYcKfE6Ws6QJ8INaBqh+RXiQF
4+8Gmcroy2lk27WTJSZrXv9eVbooMatAja2pBJsgmLNGzGPjN8vxtrxwLvXvj6VA
BC7HDPS95k9M0A/9bVfUF57+ThNBTgTPUUc2/iZ1AJugkW7qZdVflZEcN/zAn4Hv
Ad/hLTbXMyXvMXW8Muj00vgp1KJMgX13g7YDDH1FAI7Tr13jtmXz2qBy/5tjZf8Y
TSaPadZSFC3PNU5pKvTDva+2Ogq5k/70ztbuJ6B4z/hvVtGkDLKE6XAvorDKb1fq
L+ub4CdpWmHP20muPT4bgliNefE+SlegXyrnp0NOT+8w+oaHUtwvGsGDSxc11TRA
72YP0rY6t+gSGGKYT++CQdrTP8KFMtnJ814z6DdE1PgfWC+6I1ciqkwaVfclZ0d1
dutrdGNpmZ5kkB5DCkere7KikgXlTL9JNRiU6e/IndmGQNf5atvKxzVjNGp3wwPZ
k7dR8F7YQMHOCOecBjidxyk/ldNAUWrGq734Xxpbdesf85eD2DjHzJ8zdlv1Q6lD
kmRWhhpBJEaCC38GnevqlONT6AP0W/M7XyL8xxsYq1RpjhXL+uxAqztnLfLdtH9N
T4rt1f38EtZbjRkW+Jj2FEUukCkLhwd4wI/2DEBBqELFvCXEvlnNPxCSbqG3VjZW
Uaf28bW8b+qsXRB7Pto8flL46JsbxW4vD4PF551eojJQxvRzAlnGf8veHpf76CXP
SU8BNVKF4Hopa9XO+rl0aHQlKMvPeJyRCOf167kLIBAuzIZjgmnPZ24WGzRqtolJ
kPz0nJfo+zS6jP9qvog/5o0GKebbZt15OjkeB4fYyRXvwAUAtqivUVewDfycMvrH
K8BooaQY2abAjxsnVyRVubLr5YYT7N3NfBRIOg8hz6RcPMIlIo286bTs5wA6s3+Z
/NZyQk+uYVU1tLn4kh/UIU51snhPUEXjLduu8wIwpVFRybzijPuDrrKEhBzf1X5y
1N1dzWAPTYeATfru1lrDu3bblD25/JiS9N00JSSRhL+8y/E8KvUtwAkGD+au7YAT
E3IkZzNgEaJ5nRGd7PYfhYZ+teDXcrY1XJdv49je+w05DAl4Bs146SUecvGgbrXa
00x1nXQdw51rzo7TykTAkdCgfxNFs4I6EZY50j2aKBBTQvnTuBxshqR2rRNHhAgs
WGTRrEiZcp2+d0N6Oer3IPKKzQZ0eEAGqt2BboZf+1qZebFeEJDUbJrwlJwMVtfz
gcRm26ddRFTWZxKlHS38ctPcbqu6Ut3QpodAI/LcJOk6n+brW+/EuP5STIVLSmpi
PTlNetkADbObQ3bzW96w6dQMjOHYsYb+eeZP+M7siPXtojGoO//F5uQuvp2cRmQU
EmZnS7cV0m2lTn6Fg7HueVMyduO7XPX8T4gHNBJ7v8tL2Zk3AbOdxxQXaBAm4lXf
EXnVgmKlndZSfoQkEk1dcU0ayfny+jzC1q3K9y0DGVcCYQW74DRsHYNC8/33BE8C
hM4RfvaZsv3v2WK387toVlbKhMKXeBzWXLzz5E/BTArNTl0bB38y3X027JN9Pgfu
139zzyxKPhp6hSlrgCiHBP8anMrcxPxm4fZvrGi40q47hCRpCY/FazhayXhbkY1Q
nWoLhiM3E2ALi9RHAL+QN7vAvv9zwdjIdfgdYg8PS9DbdeLc1j+55ukoyOtTbsZ/
ukPz9870cL7ngdAGJm8jx0a8CvbjLglMrM0/t+aMI7ZuobZgPB6vycxPS1G4Ovzy
BRjavq1+csYiNReEn/LSum9Fi9Vrzsn7zLBr2KrtQQydMoKMWjWTM6/nX/4qWE/C
6DzvxdSh7SrqNv3qZ+Qgfoy6F0I90x9iqpPTjzZCxKwwlJfaAX/k63MPZDyQIbTR
uzeFRfvTj2vJUCEKqywCRbE5eO78zV8toxLcVmN9mQjhGxUubvcmDq3fy5cedLI2
ogC/CAPhU0IQlQDILw4hdY7f8CX2O4NIMhfACwgZcqCTFhEaixjpdX3XT9dZvROb
Lc/4jHCjo/SuwR+krtJir/sI23ukTqtLhYptanjo2pndsVzrRMR87j0S/77kqmSp
6fYWtw2Hl2YywJ7zOEPgCPJtziy4wypBNaFElq3KXMASbxqpsfjWSg+QsY44Ivka
V1LkdirquFYV8MI6G2vD4DBj6FG3XxNVR1zOgZUxbgIBQg2KPCKQ/exmoAtORgmg
1TJQCi9cCUCUEch1NUBlYgVM9twG2EnWqepqww1pNjOEgHsVcm7eNS7A4x88z6yJ
rNJ/P1FguRE5YaWHtMDFpUuoWyCYNx+AweKkIXaOg7SlhuSaqmfhdaWD+KJ7l3AQ
kx/l0n3WwlT6PucwDAn7huOu7HZvIKkydWQYJ3URZ+QPUA2ANEbPVsXtZwY227ad
STwaL8zGINoXzp2+v17ywShiGzoFb/70KE+fR/xgegzeyW9jNM/juhJ/mbOtFtjZ
x6PFrMydBGxLVlGfN/rnF2h4YfIGe29TesCGT3n9I2KnQjux/VdA0G0i6erj6ZkW
0na+8dfblMq+RVgfsnoDYMET22TdOOG9XPQHfCvTI4JM0TIGW3jB1DSoT7FipkqB
eW/GoJop/bOpADr6Ein3Jij0/j4E2QrE6MiSiII+SJ4aexaSd4AwA6z7ykf1Po9e
mIvWzvXGNx75EJwcBkd7Tr7vodzF6i3j3wumpsJblIP4QucML3jL0c26xCUmPnCw
1knqT1Uvcyj7YoavTB8P6KqmdJFoSShQsiv8wUO9nFyhKl9rsg/1FQN0u9x9tn3D
nWOSaidUGOUxgR82UntOqlGmDNTxokIltJwgfp52Fdinzi4V1FKwD6Cmn25VYMPq
43LEurNrLSTJ8tsyiTFca1OkYu/Jh8Ic/LTREeUfZHbJpxFBhunLRmECBoX0oXDi
Tvwf+LcxO56eTEsIxcfqxyxkR7H2+N3hNNNWYlsoAlWc4WDcL0xCMp7/reTMg9+V
KeuymywPVkv3Bgsbepz3YsHov4vJfO0R6jgWXC5RGT/SVlF/G3ADDWZAUmuNiKA0
p6cZ6YGunK2PhahqFt7Rr7VBMyH5O8HIuglZrFMT66jRwULVoRMWy33t9jdrqeC/
ZQmJiDhqAOHruBJ9AIwPyEvQLwd6JJcwFkT3/xUlaF+Nw7fUiT3nn+1Tb+cfUQ0F
lV03cxwgruzi1gEb4xZZG9PGNrWxAOQvP6rYenCLKAJe+aGZxwQGVJdXLvU0zGDI
8C8Xy2ElP9IJEGpFpfwp1RydSt9KP98ZPKnGRFRHbiSyEqBiVyrfxOc8BHF8npjB
gvbxAtltIbv1rzxEc6u9JgZG9rjm8SFK8T9JHuEqmy2uYHM0ShfslsV7Wc9z/nn3
iXgODrpHi2wBmKlRX3ga3S4aZx6YIozLxqXlP6qXp9NPVyP0FpxnP5B6m1iQ8RxE
nXtyJWTD1qaVsDjWMHtWwvzxak7cLhpmfynpNK2tDXZizr6kVkDPVNx6gOGQj3vP
Jb3dHz6qdafo0Mg9q1nRF/D9XLcSE+Yl54iDRlOWpu+Wnjxj7kTRzsN/cHFG7Eqt
PImC0lMdmBGaDzfUsv1Ec+m12y8NF3gmbX0ShprUACMXYRkrcX+dHKQYcOlK2Wog
nCz2q5VLpD9j0YrBJ9rXI/XYFbo6UKEsvQosjb0v9cETwn83dGpRqU4lrJetJG4p
lIThf9aHRxaXpU1sswWhDl4zlV9i5794+2s5iJq80+Ev9o6QR0TMX2PIk7aL2E/0
Y8Ji0K3Y5Pt9/KCCYTPdDBiSrzeRum/AO1G3DaOJQF1tjdf2uAjdhIzMrs4SpWyf
NBVuzRHbMfsIMyVocBs2sZuvsaNSYb5UxUxZUsM3PvsRtmdHP0I60LqgyNDV47LQ
gjHYFI+bthKR3yqIo5Y4mimAW+Vs1+VgDYnWU4rvw3kIoNpiMF8vHIrCiMc4sGKW
HqVYBqP0q3S1iYuYuVfKdCV+ixrUGOHxt7YxSDJhSRdmNddyFixTX8rEgL4k1NWj
UCSM66As84tXccACeUm2RNmQv9A6FnA6UboVlDBpALYbwxw0pZVnK2bJz2WYs6N6
L/dQYQRhCz/BKhLCy5YSKh/WDOaO+YfImrcpnP8wo7eApccQHWREQhn7BPXtxle0
MzBgyjiCX29G5dOI1rShzs9h9jSKDyx8wUjrqwMrA1/3M9fYYst9E+Ze3amH9ZgS
FruR+6KhzJ7XbNmd7kNCu3O/nW8xho9+ZRJTq7RG0lVcH4n5gpywiXaZuaTrtbMS
hFutrw8/50iwEQZc1MsadkvEkWEctkO/J7Y1UfRaGTDL+STicrMtl7TS7kA4zn03
+mAbWbvYtC3hJFS5+ycB9WRZmoYem/cp1KNYAzdxN3s+raeBwadtXyGBMC/3bb2c
TZFKO4JBiYXWg21PmSb2pIpByzq/Lnmt0Aoam3iTq6UYKgXioC5tcP7sBE4FIh4F
VnwhmwyvQZI+SirLFSJdc55xSlBV2Eovx2rbS3h4RNPhxZfN4CmhmuMhG36b10O9
LW87ItL9Az6so8mUyjQhH10oMl0SWz+cO34l8n0HRMdYOEY48b5Y8ht0ZKo24pnB
hnawA9uAwbBaqk8Rw13x+vgS6OvEEoa5pWZZuBqc5XyuLuNLd9YHV34mPcIWRmhe
s/hro/HXfuC3gRK81821JtrOjh96dby5ExDJsiWH256M5CS9koifXWHGRPfqKqCm
ZNYEFjgMqSB9r0nmiSJqdb1+7n5oynAmGnSVjlDCtLcgZb4lpv3DmoH6CN1OLlmW
TGxY1WmnmWXqFIKsBCskb+1KcZu4hloCGphSM1A06jMH2vgOwuSd4liilo5UqjFg
Tc4T4tGtR8Pjrt6sUpxTJkDlnM9ysdTS0VC/bof1X02w8wBz7wzeGFJUKcIvk8nt
g7iRARA41dK7k+3hsrtLYf03D8/+W8rP1mQByouX0Lr6oQ8R5ntZDW583Gr5LGzU
H2pbuxdL81qgDu1ojSZxdsmeoihSTrzb46Lp5xwdjpAI6TWTmFoZUCnUNcbQvBbW
pPPOFcLlRHB0DtL3MrR7zWbQptLi7aQoWiLD1dPx3gvLo+95rjjIIQAjnQJgp87S
2+Ft8++UH6r27iIab/NtVmxZQfFeimwb4wp0z1LYjUbz0GTI8OSdGClMorlS8UWJ
z23nY73tdHOQmJd3s7Xhg2NutKpL82P/5rB6rKtNd34DZ4pZHwTKepUY+KzZ/etJ
KUg1d64EoFQ20TtJJj9AMyoaZuMawaG3W6y9txE/34YwhcgKVmxLkL8nfaYZDlan
Z4YwXV4Tq8jz54N3xazxLeIrhHv3vSNaAqDNNlNTHRq7anpoYI9x2CeeepgdmW64
ml62K0017IUtv+Xa4cQlnK+dwqLkNEjaMGOtYM85uaSnIewGANUevZnVGaLUqiqu
OHsOSVCmjRWZpsyrqRiVn+XFX79sSwZOJjjdowJH0DLVB+DpOFbB7XHZ31N3nHNG
z9hdJlig2ePWINZnx5pU2G+/mNdk+cMM0QNKe0kDhGvEgj9f9/oAYwew3MzzDA9I
fbBf4dSfX4MhH1ByPuX61aE5uFHu829pisw2U3IEh4EkeSnvQP/wO1EYrlKrmK5k
XYRxzsm/WpVPY99ioPJB8ELwxnv+/XitHgcOfeJLNQW5Av2zqjxxwgjfwgfTnj+9
aLZt+0NoxKMV8pGn/BYgCMpEdOdqHR9EzfuCT2rxPvg0UGc2OviyKT4LxTeb1E8A
AYkqRp3dIhkbbYczBxqkRjDDUdTS2I4NAdL1lBV8uSQ2EX+uXx0gJZXCQ+h32hly
aI0vdtknnHye4EG5l5omsBhjIJxJJ7h4+THxeHX+i5M/xuikuJQny16t4EoKA7mQ
fsmC4K7OSZHIkyFY2Rsg/sNQ0b3UUa/TvTUriiZ81KXnqKa5vPyl9t3MROsbIiYr
FQchEfbv41m2Z8Hda1tsnozbYVxdtxE85ZN4BIzchuHMo9+qt5xzfu0tCejaq3JN
9hQ7FhHCZg+G940lpci0nN/8YYUImuVNVSa2AxFcr6i+gLiB99QqWNmuZeRUtNft
l46da11IASmVbzmKvXCHn1/mNbXyMeCa7u7QdCqUI7+t8OKtAkbXGT1ZdiTJJv2d
ZlPNSKeX007Up1iF29tPossxE0uG9L1BC+sTK930cMga0fmdy2oV/cPxPUEYoZ0X
MpopmmXuzrIEZrVNUBPYUCHJJDfML5mhI/tuVpYBP/yhIMxDo01WT5hcOYNWNXrA
iYnWY31uglBrKLj72kyeVngEM5BksapaLoz3w5baxXjkxAayVvbRgLT8ev/WUIpb
pFi6b53shRjl9KkEZ8W2cIrP5abLzjTTypOu3HnSqbF4TLlmXW0q6bKMK8yPyKox
kuBgUsL7z9xjwzbcWQwXqwxy0jEfAdLFsGSEf2Yd1EwR/ooCeMmRPpFbhprSXpwY
WdokahCYzh08tCxEouQb4JXcRPYzkz9+zeqqW0WGHnIZP0N4JRBHJ/6bE1ZOTjRv
eJrEo6iXEIY0GC848274J4ixPoBH320Hok+aWayXfAq+IWyzzqIoPek2KB/8fP3U
DcVv1P+CMRooJj8ynoWyueapDJj1i25RdeOd+7BLD3ADX6Pbj9RIM8SRkWpHEn0e
qEmz0UTgct+TXoIzor5NL1ins8zBi9vxxtaL8reiLi8sFsB1+/UD9/YbZxLRRYJd
cUA9qpXYuLGpKzXFc7KleQgUuK1no+yfvE02aQogfYTi6PcDCf3AX9rTxOBPa0Nz
sOA6CTlpNjjQZ3hO+aG9unj87P9AT4scY36gsLnkzThfRxcIaYVt2nDs14uehZf2
mOHyhEk8O76W2BfpBRqXTtz+jR+ZmypAaEZ31nUmfTQEZ8hUgslyhrdEOY55SFxe
gI9YZ1CFW3f5IJbQvwgrmKmTgxr4lhuUgnsRHk3ELXHE5q1KWjMUbXCD29Mv8hp8
t2eKBMGV3310dTWmIB9X29mQ8nW1lc2i/mZVNeIOLRymdvuY4qWDgXBvQ9C0cZG6
prw5gcvptcDcRj6z+DFkkb5gltCm7HEcdsnf+FAb/oNtMjCJM62cTBX7IIbqcMD4
g+/jOLAjIzZ5H6LJl5TT6XwnHXB73DnXiRsOvq0yKLV9XA4k1Lqw7V63b/jY1mE1
jCE7bBy3ObkZ3GVEkfov1ik2+uN9Fxjy2jhA4GYYqhGvJB73ockuuaNHY4pAKOT9
IEkkPVlGUvTQ8MsU7gmT61J9KZ/Qyn6ENGfRWXpqkS3mdwjtrD4s9S/3HbcEcbZX
TjV1vjoEFl8o0EQZQdrtlLvXi7i+2SCdycLVJyb8YE/OwyZoItbClqTbXI2DiFhX
3vchsIXNApirrEa6LX4r1FUXxrDWYlCQMoeIZnqOMaKZzheWWIX6o/njG3omhCIc
wRC6N97uqsRVaep/KifEoe1+mf8o0FlXD+XhDNomBtHwMPO5xOLeb8So8iqWlnfs
3WSEUyVu4Y5zM3Y+iMg8KRGwxiYB61mnbhP10U4e/LVXPtQGDHQzfvU720JmcLtW
pVtiycrhZeZ+q7aFU5UnyIHxjHznKgz7THxO72jqv11JBnW0ZrqC6x4XJZYvDwst
79j+79Gq0il3d7nhIjOhl/1eUM4dMBkU6fVZnUqIgU6RKhtNfqNOVLZsWBZGaOrK
hlXMHaICgbzOHQa1CcKMaD2XqYdC+eCj+n9+SybKENNugfVx26GTfeI5SO+pa4UT
uxeoJSVgHvgsPXIFga7jIklMfcbj6LArSXabkW8tYC29XaG27E3g1ps+2CEZMHhJ
fNU1a5mOE9l/th4goC+/ZdSgDz7rNv0gI9bV+s3u68+4qd2TMeNqQOWOEcMzID82
hErRp06KPlSeC6P2UehjcvnUbH9V8StmCf40OyB4z+l143FPAAMx3dThy5tDIP4j
LcmMLxKlZtfGNoGtxnCIYLu2lkLwWAIV1IN5VO0pLufZppRWyyMdmxqBfYKXJxNH
RASCbLIWdJpHOFIYUUvBs3lx8x9/TLS42/Tc3CFDpR2BCsWGtretazssrrAVX4Jn
2GAngZtZsFIoAG0cJC5sj8fbw1gA7Bp+PCPJ9gOYmUTylELBqVoJqj4IgX0LBjn5
8vTg8OvQA5VynPpn68aW2d2eaY7LBo8hFviAg5TbjTVEU4YSXfEM0gVoVs7sMg1U
7KQIBjPRgIQy1b7Z1qtPpU8Kk4GhOgmumiYVieGMFw4ChhZBcOvLD28EdbGO7M/W
m6y83XyvzswVwxt3n0Ke7RgaYyFjXdemnoU07d3IWr7kzJEXcOtqbjSOVZ7vYJfw
Ahh3tgqW2/jid+lhWuvhjydCUsjWQFl30h8B4a9rvV8He6ZSeuY/MSRnZcVUrDwm
XJjO9x0EMZsDFpg65hA1A+lpDa51xMp/RP9YbW3+zSZ0Av9U7gaoGXIOFQ/KQ1j2
6ipekjiMvUVn4k0ay9ak0gTkQ+wyJz9pczQN17gU0KnS2DhFE88JCo1bhhS2bJl8
U7FoMip2FTsy3lN3yhdXpTWzMSoiUa7xqPpYufLGtQVjEYnVLItfFDig4RMLg8C8
OG1qiuZosixvMqyzHnLxs/iL8yVAvvoSA7whaVZl5vxOeg6S8mPxGOJaqIepr+1P
bop0XLRgwNpW4Ggntqy8KqHUPPVxMeIqI7lKPi+XXM1mndGZe0sgmu73lhFobSL9
eBSzEI3dlUy1f3K5QrTOuQacJs0czRxS4dgZn1Cl4AJ45/HUZ6xG/TOmauW7cVof
wCWhVjXlRCTlcw68bi+Nf9cYkHdBdwosT4JHA7KZTU10QLYpv3WKzBZ0beXXVyjQ
Iv4iMsvt0QhNMlYJG70q1Qg6YBVXELGePkdQbljUz9+oFnkQYR7o4SfuI/+r+s7k
ZeJ8QfxX7fFdnv+4maPkwU3PRar+8MUoJ1t+QrBOtvATo4muAxVBM7uTZWB+0UEV
lvKbhjM6ejxC+9qdGmhlMF+gVIY+0YWM5UNw/F4mqo1H2VdAAmx6xQGQV1jdko+y
3RdmyYxd+qbdz/OrPxL4g+mVUmHTAXPGacMsrDDKuvY1u0GIlDHWdSVfDMs+HhbF
aI/548LdfwKueRWO2SctQ1+v+6Xi5DP8N33vUbLVxpKY4RxXQ050EbsWagbA1/Uv
1ntztZXHukGW+L2ZDqGI1kbUFMjW8u0gmpBjJXZe/agySBJE6TajyLffT0JA1oMH
NYH/4uVcsPMN//sAN9WzIDKjsh3qcqXnE5jCxT4A6/+WsjpQNw06Y+qVRYDacanj
XLgJdoNmQdjbyuzMmDwfTfi1BLzVxNxyrUOfhbEZ7A5+qDhWzTf/S1KpRng5R/f9
2FYevQ4FiMzfZKJmHdKR4EwHR7Vu5YJ8FlDgX2rvS1IG/CVywGrUyEsd9hu8MUN1
6W+rgYpsBwP6XkI64X2u0fNuj+IlI6PXCq1gXrwcDqsyYC8EfDxs1ZbbQgxXifW6
Re9FiPEK9Lq3a0YJXYlNdOq0E8w/F6jPYniaaUmsc0ltQb6Z8NkEUssnKuZ4BHUd
fPvNhJWFBrHvERB9eelgT8U2GFcBw/68gWcKBLmM/67Llyo/K7ZvNTJ1DLsYFklQ
m5/mfmjLQEc0I9pMFoNHtGiuPdJigaOjR9dcNybB14cNr6hQl/zprVk8fUAT11kh
2T5+KXaodD64O/A5M53GjJ+Zxnp8MX3aPGoNCagL7TDWaQFoDLFT39fB5igq94wk
PsbXYzdT00DqdfUagL3OrPWrOmfmH/je8ri0c75bPZYoDmetQLcW9H4Hgg2sJMqe
26RQEstY+NgmdgQNQbE8alWqhJUT+KmRUkH1muf4sYXrwHONqfTEf21WJ/6LdApx
UMMI114mKZYFa759zSKx6dPnZJmRY835cs7JqlAWWB0QpxqIjnxnKGmLKmowvIYq
OzReG92UWOwkiEI4uapOiAjtD3MtYu9YOek1MHk2RhB/tvY7wqo/oWZJuvF0Xbjg
N5IQgQICPUcc0DbFLS6+R02dX7Jn3VhFtaz5NOfk+sAznopJYBY59TfbLzZxKx5v
Qeb0dQfSExhFvc+TYQ6PM/JDhSGbQTCOqTsmZgsp9+E9qKwLWLs/lp3BjHOAfaec
lNis4deVTadZmtRgdzslr3YIR0zouvuUwSsVLioySvjbhCsWP8Mu1JzlhOD5n/5q
/C9GY12ahJ9pFg4ObsEhADyc328nHCd7eWN1jcPFivoSiT2YKT1oSPxq3nOnCSEW
WI69SuD0qFduDENg2hn0gSNNOEfbLgze7lpVB7LgQBEn/XDGJHTaEnNiEwgwuvWV
ePx6EBk1MJ5QiHm1VudwgM9v5NboYPG73QJ+QJCg0hOUGrmFRmctWbirovdlr4x2
aTk+YNHnnK8jpPh/D9z/jox5Y/msQjKvGJCWnv5kDIAU6y1hF3PDNhcB2OA5PpVv
PHLOs9ftD2OyE8NUOKP1+v8W6LQF9In/z8Etdn5YW0VN5uXuWzxt4HrvFoSgThgi
PYL3p15QC+8u/y68++xskofL7Rec/R/r66f00iBJwe5zaxbjcJ49boTnZ8T4j/l+
tlaTrTiwJw1t1Ln94vfO2xTOfYEIBTxbXkYrZOJlmE7FBpsA281tBjJUSiOaJQDp
IbYqNyWlRXCVQJJSAlTBast8fJ3Ug4sWEGwCmVa7rKSdXUwNdvtT7eZ0M2avAebc
LCRRyaRJYsAOa8HG3fWgFJ64sX8/sQLSKZNFs30AHHUdLJH32HoL+4XB2g9YBpqW
uexWWXOESv+UmJTK32G1xgDR2xE48oZ1WL9WrFEsD8L2zXcC13M26aSdPmR7S9ok
74blQWI9TAvsR4/n8h/xUr3InLHG2xKBVqUXKAnwBtodOvjBjgXpUWQ7I4/naJkq
3Bf/Cl72R9o4zC/GHIriZOVLptv6CyUSPvpie81PPIJ+Yxz4/LjA7Zc5LUJi1l3e
XRikyFS3V8XFgUjpNdn1ZhnYot3QR2U9RwqGpK67katRG/DovADeAag0l5ZvH3sT
2/w3NUlh+AYzY6S61Zl6v0xZvu2sDEOdwe7yY7/S9qKKl25RB675Bqd2B9AYdk8T
IrGRY3qKZ81kcxIS+ZuLzzD4Jofxm5E3gj4X+P2TQPyctE5OhVWrVs0BtwiaH2QZ
eq4z4rIHBDVRezTaR9sb4uQwVi1UNYfCPwXGm4kac387rrxgvCvpMU0l058r8OM0
ziiRwaN2KVPuJnqBTuXG/ur5+9HkmRfT/HQco9mcL0AwcaXyVF9LNd/5VeKEHR9v
xYPdxHZeVcsE+6GOWIH8k5DGn2NzEhlBFfqYPWzyDpSMmWJmzqYnS6lfKG1FMgLp
KRmqDmCGMLtnkowBRt+pRMxGcMxZ6tpxH711lZ46aSZRy/PIvCFinvRcb41J7cpr
F7dySd9xGzqSm0w01GshEUHz5rTS7u4I/f18FUadV0tNeJQR1UXZ2xoksT6uJ7uk
IvkTlIpMDEFpqxjQmbFtVVLA4qwslun64uer3tNrBjg+CvH2nDRuRSEVG3pawT1B
2+znYz0brKvHU4jKpRkqasAOrqRrdTRaSMg0so3+kiCBdKNYUf2z1q34zPoW7Me3
tWvL+iEsSn61q5Z49mRPN4GlvDcflbHHcugPwIYOyndUcaLDVBAhlyKQ5ga47qeW
MXcbbWCsjJnd32uVW0P6/GqmdOieowbmk9rs5hgUBboXviV24VPq/48kikEjied3
9CkiC+xUimQ0YnGHSiU1tenfNi89ffPn2VC3hXgLOHvHBSKPH08fKptgNvQiL4IR
QRSpwIkHTG0ozts1IGgTeegrwWiKTl3jqD9NRQrm8RmoP0oVuUVjffBmZWndPKYh
2CSG2ZX2J85vgqXH9W4sN7PQYlIegRrMxv1BlG3mnwGj0s9hb8YR1zvrHXwH0Ety
Mre17gqm+iDLSGs+pzQuIkOVu4dNYx5aTQLpKEkfVsk9iGxBSxXMEccbTorePcSe
qOpykrblRF6fObzip0JxVT7tFbnhnZT0a+KuszKfTGMdqtS+K2veMsVp3JbgS7F8
EB74vL2QzvqyPccH7GJZr0jAMuEAagmzKkL7Am3U98+csn28St4p+at1woF5HYLz
sJ6kRj8DJH686kV6si8fLL9VpSnmXhgjfV6R/8Y4EPQrJ2jotGx/i2ySfjiSf0Ai
Hqv7D8JwBUT6UuqSa9jYORBNJ1rXz6Y9THv7pxCOOFaL9jpQJB6uZabhLg1/UFTR
McITOrG3Yx3vbZXl3EmZNR6thzr0/I0MyrwkBDaKoCFAc5hsLCzfHKNytIiA5WVQ
AF4W4qNay6oxuACnupkeoFuj7EfTbqJq5GkVUYS6ZMkhPd2Wu5i+FRA5yn9zG/zs
MlFx2oCXhP+SLgWS7424WGiX8ytm8+SJuymzaPY3ZokHPwzb62ItHrTpercAw2NL
wFk1vhZsEZHFyNh/V1PZh6CzuUeteKkGj4AUDQKBQf9TKZ2xfkLZ3xIBa5nMuSj9
qVImoTK6do8IrVcYLKyI7FEJ2r6Y/ddxZ7CjNtHC081BHz77lui61cSQIxx9sYk7
chCLRDXXrngiNRqvkGvwsN2WT4DHgVUdRVdDeF9bsZR89tVl9ryqkfgx/AN5bJuE
f7dxoY4+XuLhpkkvrUuOYzavMVYPe+MQFL16ARY6KU6PMDjopFFXeQblJsmrNF3I
7zOUqDBjnMjFqhUvq0ia5I1/gqvg3rVi1f7M5HldIPoFEk6WQRrr8VOtBprhc7yR
sO3mlmiUhY1B3aFEHiG25/5jmr19xP9JpILHD8cBXbDj32zSjgmzFW+1nC1k7sQ1
9BHc7XgfxTU3px5T6BhThhSut1kLoV39ZY3jQW50cGOOCU5e1z1BOk9R+r6wmKRy
LGTkgXwiog9JzUXHf1gC1d6iGVMofToJM6q6xJVcJoUJD9amOBqnHiWwek3GG7RO
0C391la/7ognOlsyHm1cXCgulffHIDlis4+iNSSL8t76h/FveFOAwsPnsroeryKJ
qyxT/PBugOyw013nk0WCDND8KhWESFyUgapXilx1eDM7bqn/d00/IrkmmwTDmJPq
HgBUuSEb4+tphEtrivZIIdb9ATz8g7AjLFc6iSZkwwqRlwKN7KXDoxxpxgcvzmop
iTG9K7sshOJZyYgF9SqBb1a+F0IPUI26jUevfw83tDtoFaapyRNwNTYWfs4hpdmW
wsOjM7A6BjZqqwzGJ0LEp65P2RUi5K8NkXkHHhpSTNbkIS3618r/tD7vUEZoPAfR
MelswO7p4fZrox6gjiUZQZ6OGt/rJ2btwpjFIxg0pGGcwX7X9/klnPepGEOR9Q5J
wRoACWdOxFlnuIlaUEzQ5RirkgKZY3GwXvWRuEqISA+meOYmWLkoAwRA53XPde84
VOkgEZM0erW1kQ95WfTS2bk8bUdWvkLhIld7BxRjaLex2ZZ/Bxo7LA7YjZmbbqgx
qCPKb4ql3AI+8b2eWzGtPar6HiNY1PwRHDv/GBkKSvAlg0ALJa3xAlon2fJ+TXPn
K6SnjoK4bU7pUsHYFAOTxGzOsD4lOPi7StZ5U5a4450ZKE2fmiQeejesHzG6m8Nw
fM9N03jZ/Pi5DWkBlcF5O0i5A6zNE4TEHUO988igZ3iN/vCNncxLruVvNXlaysF4
sdJTW9tU61asyI4ml/c5VW4yjfZ4eOAKpJnqngWzDwhUjpU3zeqsZmU0s429cOMl
i2VysP/88WE4zJQfWvIOb1hV+VPMNx7VtTK9oSWywoHO6+b58rqTVTN8/AmEjJe/
yekaCua8wrGdR4tK1elg7f0QlJx76O78X24it2NxqIH7xYCCm35zt+/JxVAnouFE
fsxh2DrAY8uB3KRnc9Z3cMtt0ETtUYE1L+5Wh+fV8rLN1ob5pqnV2SdKuUlWJN3M
R8UaFtExcuaP1KUW4J1iXzbhOugkN77pm0A7oGVOIiqgcsqD0V0NdmEfByLPrjG/
62jwYIUqc2La58vjtzOGYivFHEoclb9u3cL6b5nGonJ/RCgsMO0p0Gbvd0JoS6XD
RsJkWA8KOguiX5yWdBIdSYCPdb1Ep66A9t3kY/Zb25VzH7IHqiZjH5XU4W2jayDl
UVnRyq3o5EZJLvjflU+CHqXdf4F4thnat7as1ZPGbcBUcp680ZJxMi49LdFNQMnC
NVHAQSNDiAT65wF5x1oTVNqXSWW+vgioFgzdBIjqVzBqz7c7mf7s/jQvtsN05Ub+
3C4gSpN//rx0qA5H5G7yKewp1rW5wpw6QzSzHOxmvxBOyR7heBI0rodkwRW4Ke+u
9WciayZiCusMqPvQE1/1HSDzEJOl7YsK+DIBq4JYpQPrVL6NsiM7y11MZ14uZtnT
CBMdHm5H8VJ5MsgB44NiSrGWFMuLyg1EswVnOvApSutzDvuPwUhuShNmX4liJTbM
mtAnMKdPS+bRoI907TiPNNfyMZF111nKG6JiVAiUqRWaLPpmsEHG9qzIVp9cX1qZ
o2TMB6Hux8hZewZ65j+d7D8DIL47JYi4BGsZDPcmyR0PMagnLKGgUvyiHYLQ+WUw
NSDBHcr57qNCTh+O52jK6BIl0XICy52EXg0JTub01u0tikt7rBIwGEksVAYz99nc
F+3PTRDVzPercMTYoNPwYH9GH/YKvXb4msd+rJfgSDgptcEfx9QjcWX3Xlcr9bff
TNJIF0ZjpT5/2WUEm5PSYaWsw9V1reW0iasfMwtBINFBketZ6LpFRwXB3cmk0RMn
dQ9PJYFhn3YaSHRorQuaPHo6+QGoAt81209FFTGQsRH+ezt2Jx+ahhw1RpqRtVDR
C9HV/Cs/5g69OJWjChWvIl0WMos/LdWRmpyYe244CCjiilFbG5MNQWz31wQXjR2n
Y5MSH5XU3vWo/18LgIjbGzpkbMVOb/ppHjmMLnfZL2tJBnWBrAq3jr0ppa9HWEo3
3qFv0A3DIjy0jz03cX+f4lSOkQesfBU88Zi4voiMR7geM/K1M8c5pEQZUPWC6u0t
rNQh8Ne4fcubPWx5g2MVkCRom6guAo36zG2su1LNlgetIiVkjW1kh96wMxU7wK4M
dvl0u33HwvMkwbYyOla3IK+vb5r2ZN4n/cHhY7ijh5oYyE9SR7O7/2Uzaakv7AGf
Eyce7enU3PTxFxsD9Oyi5Bn94HkOJ5vZUdTbZkrC3jiUFI3xi+Q/TSVL2LSaToop
szsPS5caWI5ZwOrW5td9zvw8659tPu+JG6gNF2iadfYad0okvGIYYOr7akdvuMGQ
4eTchSL0yrsep4xIPX8ziUdM14uQaawiPWao6nWxq/T2V9pMjDaposWrZ7pYccZ4
SQM2bh2cgyyA1I8UqI7CwbZdwbl52B1QcZaBkwaLCUKivOfujBQuxb/cvU+1+ePG
lxhTsOWzVHt/2XhmlMIiZk+79SpO0ubNYTA/avMCqK4sdzMY0G4w2CD1NaL7MVRU
QmJpOKS14bzU7tIgGywszkCGEqCf3c8/nmqU+V2T+r1agpV/Qb7yFxvXkffNoUNP
RlM7kbT/H9ee2OHgV9+n7+1uYvNejzAg+aOV1DhXnoLu0GMsPiPHmPVnsKpsGca3
zrngsUE+4l4ZD3h7BbRTdcjU3e44hkorLZBz3MFXpjYZYXbVWOmFVlHM3wMOY8oa
lZBsD68I0VrN41H71ju2wFta7104K9DtFNkixPxOVeZuRKN5lYFZMbuQWvNTgFWG
0mBejJgr8uxYWRICi2SqT/ou8VJ4MgK6WR/BVJ/Vff/JvsVfbS3RlKsHMNmwrFPn
+sC55K/umOQaK5puwMsb+6ZILALXT3lLn/iOV9GfuvZ2UEEJ2ndgz8kerOyeqVjs
apwugUkU6/8Oc43hDtyuSL8iyAIUZ8oqCCMiRbLZpbV7PMRQjRNk0LFANoFIXk1g
6LAHHOPc/Z1xXBwHdonw02b9/jYI0xHe1pDzKeICLwft1U6laLThJjhHxIky2enu
P+LLV/fNe8Ou9cTd0Am9MhZREQQ5LKBPTngD0Rq829VQcL1RUCz4CN0g7PZH0btc
/QBEDXafy3St1fshYavaDAiz9J+oNwPV8IMwdJK3ZZFah/OKcfnLvyI60kM6MPB1
lX0kLUlztKohURsdOqd5hi5LTnNQ2jow3v3fOhKftq+gwhIhMdWm5cBq9II4SSYG
VJkZ42zIjr4SQGrNy+fXgweVeTZm6iJJwc8J16AdMEeIkUllBP10sAl4/SmDOere
DQmXop3gT1x0jo6hIEZFIjR2IDqw402HfyPhLg+0zQoI2mVl11Q8W+8ZyxY2bnXf
qv9SD7rG4CJ/6pd2DuEvKRLtHeRG5G6ZaTQ8tBkr8xcMjZSfl9BsynGTwQtUvg14
JhYDa4FjXMIl+RQYPB9skTSOuDtgW2QwYHtgWa293JpAzHYzi+oOLVOrhI53A5pD
yiouBKfvLnC+U6EzhjyO2LzvyVrkk5qKamDso1q6K9Vg99wLa2vqitWkTgr9xi3Q
EB6vxS1vv6NrY9eJhMP4SyE9qprwxWE16uXWuQsAZWv7wlOsprXcalEAJGivTKYF
dRA01r1ETdjvnDGBf0TDJ/NpTWD6nDW1xe1Fgph21O2Nw0Rli5rfdGiKGpPOewLc
AVlICh56mjAT/CBymxr3Jh4A18/+ooLQCREkPeEgzSjECuvca/cNsfZI1XcOJII4
E+EOl79t/XUXc2HT+kqk81QHx2uKofguUEIWDTtm1IFUK8xlnnJ1HQipXAVEPhsK
L567iLzONGKTDeVJ6h2XFS0IqLCoRE+ptCksnjEWA7wlHM10bcjwyg+D9J6g/ggb
1vavBoLHJ8B6+DdvEVDuIriY07xmeuEXKsVv3IvDSe2/KAap6Vv/HCOuPA4qo9VJ
plgzjt7vyjewRWg8fSj5Y2qInrFSQHW+BW1R2GyoF1Tme3EYHZEVNIGd69rBCv/4
RUc/cX57N2+nc6AAtDxDiakBJyCo3a/FeNUOTJTA84NgazhR8eEQow8q36oOoTjm
56wC+TQ6kqz3pNqprzSAXqzR8OKE1qfgsEZYlLDeysiyElF9mgouUNI+ZuexEcpk
nQTxdUFmvwSEg9Pea2qArJA2gCngDJgREkAuDvQbHAUzMJG3CmoAXlyAvkPjx2qV
BRlr4LubaJctXWcgWnjFyCwvNCTd5rW4kOQk1aP5yaqSprp7ryQBvtO701YE6IJg
cCqlKgDhouIRZ/qEd2AWy1JS6Q+o3V5JCswVkMf1AIsfL+6wbC27HdlWzxEjDEYl
qKdhaBszcjshv3UV/FHV6lmf1Zz+UyAQl1UN6nJPoc+nGYD0mW0+K5g7Dx2Qf/P0
dUrx3oQOz2ltV8huL/XfRFUtAXhGDlaMgxEqrGKGlw0XXGGH7FQo2obTTns3BML3
I3p2cGdxanYmQQRDRyvR/+JhLoCkBl6Sp9x3WOYdegM7QXeQ3PkJT7NqepYyj9Vn
bIUb53Wg/pQfiOKvth6m0fEFlStXVaDhIa94Fblt9ojooiHpKvFanghceTwDpalD
PMRNBgEAO/UyGhd8wjtdSOG1TumW27aShZU0TUY88udQyqHjWFQURt2teVLBsZDt
pd2518A8VMlnRP7kfPvF3A91ptBzbGMtcQ17csBmXwzenGSsC3P48FoI09+qRdvK
ntPvRB1kH3vnqgNiGIGacFmg/gQ8KMaeX5K9QWLGbNU0hp7NR0gysyWL6lPtW1Sh
W/byrGRdBnUvg0jxtCDTWio8dxjEeUnsAC4ukduYHa/Z7pTWc8BJlCEyl141bj53
6wCOr3rP273dXdPRgwnglb3A3j47ib1sS1iLN5uVzUylxMxp8LczGrdLavOiMkXg
GwRAwsUY6eWA6ruiE2h9DGkYD4ZSOOYv27E7kHiwany437RzfLgRAFolbtGYennr
9KfGen0Ek9Y5AOR1z6IxUCMjLeGbTjYlFrdR7TZeNie9qVVehfdIid4wdXKnEehO
6UiLNm2kfAurBzEmh2qZuuXcNgXoemkitOx+lC8iFRcZdRFcuJnGr+a28JoXhnEm
iKzdNNb7Wn5skRapd/LuznsrKRPYmvjS/IkjoOTmNGDi6LxOAYlRbXI50o3ziVef
DZkrOIX+jrDgkeyEPPQRgheIbjIP9wlRi/LoaFvsAwSjNXD0K9aXTK4rWNw6fsoI
+QyOdrT4gLhRCZf/DwS0zeka/TLIl41wi3VkqLpZRPftql7b531xtV9DaTz66zEz
7JDnyvNGG+z2mwXys35Zp43tA/nA/GPd9Uex6J+PLGQoUCcx6f0XgoemGTIUo8NV
+N5+5zFx2ysNJqReQDJONRZI6S08tkzwEyKRh/SyyWA/NbQVHU3M9c83QsCZS+CG
eP8IMJTINKWqTbXlpRuymTz+AmWOq1zefcm5YTRpXOpRi+sRnByV63CUXAV/XrGI
9bhQHJU9P17EaYMJFHkjMeYeyypSQFWUp2+lzyKyDbjVDcbU3VgS0qYtaxr8rNHG
8BwJ9Nq2oLHMfpDkLibtc+cvWvJZNLn3l9g+DfiiMJ6XNfWBCCbmGgv5kd8SYhba
RnGURxLhYgLT3LOZej3D0TCa+7CtYSbdLrc46/0zLy79p350SHZOnD3UlB1qCj3j
nOLwj4KaFyaN9aa8BtqN0A7WlwK8jK4bK618tfysIHCnLiwquVr582oxwKU6g53/
0+AW/U2qLiMtBXRm0bwsrciCCeUW157X0JxYH2mR9ITqGUmKy5+oosarDviX1JvW
b3AZ2MbQXzfHI01e/+qZEBaotqjbwpfCfSaFbtFgVxw/hBFohvrmjwHO2iKZXmtM
UmNJqOv72JyZfzGwxzHgHdCqrMzHxuS+oHEzTFw0afyhKgEVbs3qKnLNhhkKoqDp
Px5r3VIx+jqYBiASmU5/LHjgU7jF/5Gb2kz3bIzRZuw12uc0ZwbD28SsNCVZHL2c
YhFHDuc+RRbwmOOxfdUqc3YwSAyHQQd5YXV0snLYnxdvridrhuM8KdpjCA4IVvnY
JYy2UVtvyiNs7WItdumQjPnTulmLnShdZ0FTAiTJHuuCDL6TaEdRsJqelbuuoYYU
BhnAboJTHRhcTXIO0nAHxUV5dqRVpC8Xszhdqgj5MAXUCIQu2LIz+QJskHu+AteC
Yut8CXo8MB//YLwp3dlMbqUdBqCVPGsZkhuGQpb7D8iyx2GLrx7Lft0msClS50G/
ujy0YM9uSEzXXPAafq7HLPkZIfGBQ8kQKrHkcCGpfjSShCEfqgizO4EfMAYhj9eK
e0lsxwQpDcP09XGLyMwq351N4vU3aaAWwA/jsH6RZoWOb2a8wX48Gv6Vt0PEXz3w
0B5Xf1HfokITMFH3iC4xTfLx2NiJicR/nvZ3hr6u+J4VjLmh/wdtfKPIzTXBH24R
mQEUtBuDN9X9TerFqEJ4x2j1xbBVoGB5X44LSdEw6q/I61WWOk8s6V28Lv6PFl8p
1icYOW56DGFvQUuN+6WDPpggGB4lrbKNuZ+LiVasZYT01Uva0MRlsoOyQteDzMH5
1kKOppeBo7u931ga6iecsM5y8rF+HCxTHGGx/KRmlqsma0Auo4EJj3+h4BwhPvxS
XUhe5ORFJFjCVzqwpSPtCL3cXwu50qkHCbFiGgD8S+aem8mxnFyxsHuK76JWQ0xG
yFrh4TqScP2x1HG5BnjyvFovzKEWjJMc/Q6yz04r79fNjB7pakoysLz3tX3gahQv
mOVrD8aydrQXiSYQYgmBzQmi09P32mYHTniQ2GbrOIh/BIEUkCaAuP/NwD+l34ld
YZuOSdhN+9lhWCFHICowyAcQxlaxh/S1owFR9emDb1d2ACoqR6iQJ4OBZhPYEHLQ
FtQ6pDeF7rSzslwEmaO9z0bjC3+urI6MP3uZTs0IYpNYQ0tGx7Wy1LRA79RuZ1xt
R6HbLbZBITigUGfeBxUoxlGDzfScPz1VCUpe7jO8oFajiPOXdNy7um7DVTDU1QDm
4SxL4ZjTmmhVvWS4PAxmHNh7CEnngxLV3l0g9JAOH7a8P/CWY2MFAGNsXV9IpvJl
tn+8WJrB6rmfaQBgjYywON+fajbx+cFjCyk7ttn47rIpV6Tte+lxYggN+8rJt8YX
9Ej9kmo4usLg0GycLxYnlNx+cyzUQv87egI4uBoCzd5p+tls/I4B7M6x59OK1MX3
6aht4Fv3AVrTiGml1u8rZaVPMzmXFwKo67xGP3bSdzvJCTvVesGPZrwoCZ4jdomC
Mj3EneCd1wWZQZMP5HDcx3szkbam9m0oTk/VTsY19cXbn+pyanfJdR3+4UlwOxcZ
8dZv4aWCpoJ+yDyd5ahPq0FnHZmlXuTAPDncEGeAHl4YYln2a2/2WDmo38EDA1u9
b97q0iQ01nPY2z6H9Fbn9oQHqzWHesTSioZeieL4KfUms935XyACGj93rFj/2eGz
SndqORd3xWr4Lo98H7cWcLiIJ0v/guDwazWDwoHBBbF5/+kwAMEmIM7igvsJ4i/T
vcSNtB4Z7S1HR8RWAHfr2YzFWM4KPSKxlPQ/0G846S6Y1wiRf4PnHLz+Qw5wpwhS
CpBwQZwxRFVoL3P4dpff3bYkOcGIw1J8kYBWegrKGgEa4wos6uJUTvwpzzTTW60a
gnOWOXxanKkYgkhIvNsygjMx+XZiUNne5f4bMvrZZyqjqkAhLlm9/uailsn2kkFy
BfPzSobO3ECOjHO8tFF5+AAn2QgfIVZJwjrTpsOmIRPkM1d5qBit8duGp7xl06nQ
arHb712QrJ3EeeRZrkIHQmB0LECZI0R+9MiTMU3CN5d6SJDy07ICZ2bAGg+6J9Rl
9EE5tjonYAXIMWM/R/wT9YRJ8UXRuBcev3opCYjIV57F6RReuRc3z9Re9LudMJkL
mtbBoTOjC7Iwor2gnZPMFzNPMLBQdFy2SdbFgcTDS5BTsUIycbLdnlKx7OzBE8pd
3YceY9+7FMAr2C49e0MqKSCgI8RqR+Kkg4wOyG8d85/Yovk2jPW8ht9IDfbnBBfQ
EV2rIeRvvoZheYJJzFdSaBIYwgFoLm3AcFdyT8Upr6XObbM0/Q0rRMcIScg/cmD+
kHz0lF9pkQ90OcWGPA9lmt5+paIzXmF8je9MclwGY012eSjNZJe5NtdO7528agIx
HXWPLzyy6PC5I66tKMxNMNc4bhKMOgKbyk7WlnD8jyzWB2TxCUfnG8AChB4pjWUh
9JaGfKupU51Qc9by37hwR3ZFHIxt5Sau2ga8JJulf46c0DTAyL0dG+Q6k7lLLGJo
kYy96OQAAGl1gd3HcZVMgwl0jWJFtTNF6KK1pK5KyOB6oD7J0wibXNLmztRyTuXI
2KKx7Q8P/fnJS5pq53B7kmAw0UYLGMJRi0BGi0h7sXjA46igIzryWSmNB0TpC08S
KB/1hD+D3Bom9PvmdJKYI9wqA3KTBTL69kGHciok+X+kDEuaLDmFsJHIBC7Z2aF7
D2tRj2VhFEYeX4wojR6N6uFk0XmH0GDlhLS0/x2rvoBbVYtA0XrO71fe/4Nfdedu
fsa1l8DtkmYLrtK7YAzVsTdhpHDOyR2Czv4S1eM1dERV4ZTrBzg0czWu8oOJN5cr
OHEfGVZpMNMEHh0mVbphmskDIDNRcQ5XE7tErH41S8NPJdKl5c5nNkbr6NqLTGJj
XSl6Mqoftka7wRCinQQqItxQsmKRSX+P+m4h6+gMFP9T0kK8Skem+fosGeFuyj4Z
AQgB5Ay7PYQNME3J5btQVyIpyGBvEIIjN9CLg5r+NSJr4/ONqVCc/6JlRgJ7Mdgd
SmwlKrWxtgq1CvsazKZz6QNnvx03Kz8NCxkgn6DLob+CDUIj6wuCDztTMucuuYjL
xG/45gFG4UjGiVkt3BTnS1PNIadMYB6HhemRR+RKb0l1WUzCoJT15UhBsMP4Ucbo
PmDR8jLPaY6eN4srfyn/zhkZHU/TFgIHoT9G/bM9k9rDm89a/Jc7jNMhX44R0li1
iPHLWpdf8jp0bxO2M8EhgFk3T9AQhb85lBxqASRR1ni0xTOHjN/Z4pe6lUg0x4rn
aczy4vTeHKlOu8CPhesOrKQTamh19YW7rzY8vPJ5DnVUEaG0gHTB1ZeIcQhokRJr
YpB05GzD2aDZ8OIHQIJijqzW/15rRYPCfEm13G/97Oo2rq5i2RgRRw3A3Pmpm2g5
Fzid4JT9I0ic709qO4oYtYu2iGqM2ye/n14LO6J6s5XqEZvnFcy1rgA9Iszct6Tt
mZQDImaPXOTULKVYc9MKre126LJB2+nlO9MuZIOY9jrybkq4GZZdn3+es8ImaRTz
pAqFBvaWKUUGl9BfI0Ol8CLjgl0fP9l1KAaKiJgHqH4E+2Ngp/9RrLvs60jhFuzA
ZxlcAKNuPuYBoeJp0HNbYEwarMco14Zf/YVGUt4ndKDVf36NSxRK/m63Xv4ddvCd
P2H/BJhsOtyGKUcF/9tT+9CHmCzSocaXTt8qvPZ9c+mdEgSf1hoaMOsnIG8XqXOH
h1een/J4rqa5OiSUPZeyzEuhPnFzQiLD2J4skz8ja52a3vH/D44bPB5/JPtJBvx8
euj1MWdbEQO9w0Vxw4rXpXfK+nJOcGFwZtQxBfcBCYbvyj9d+Bf0QyThTrOmInJz
nIJ/bMyaBqzyT9Bkttv5f7x9UVn4Vc74Z8Wlp996rZkPpYMTrzvn1pxFz5/gIh8c
8SwURQSNfvRN4oiw6j9bramAAJ5M1S9HSEhnZ1KA+IUYuAb5R4wMRJxYV+ru9TPL
GwY6zMSbjAzLqfSb5+EYJ2Lsri30ZVx9FQO7c1FzR22UJjdDJSZFzWkt6qxZVOPN
iVTTTDBYq+0v3QubaLcmc400orZdeQTVi6oFFiyZnQxLEeeYAdlANFTCOokbbitl
XNM9A6vJSGUo1vzpPsTy1jjG8VquCINg/qFUjs0AgRb+uTdHJ7DC8xRn4eE/VPz7
fuB+fOxXZujn7Zcw1TaoCD9GJUMEdAmdmRJ3su0gB0H5RsYRRBk/GMnxRKTC1m+F
j2rosF9nxk4AMH7jcNsPI5Pt/wSAmGwiB23uhMmicfYYqmdQHAt7TLISBGO6cls+
aWNuNSyTt/MI+Qx7Th+4E9l2HKr/ZZQKTOOc6DGuSuD8K2T5kIJQy3DVbF5q8m7Y
PW9BOp7nNS32q3gPsgtsHxnAMpNpE5WS/j3ysXMSbjzfbuOZexbCUpt13CPFQZDx
nACej7ZtjzI6X+K0Nq+rpF7+gU58gIqFDyIk9FfPlENLtz05eV2anGQGk0f5iGov
FeICNA5JINMKu07sYlJCIUKvd12FwKTE7BJ3ON1qA7tr/yqa88WlUHDXLc8rED5e
HzMG2ApXn+RcfvJlnyjdBvBCrSSafo4ByqqCum8xc7XW/80VpsL0DCmGq9gP2AfK
xmWR1lsxbsbqIu+9v7lGTuorGFFxVoVYbcvvVYyJM2zxOrzMbBXzGSMliOPq7Th0
thyzslcIJ7Uzbnh3JqLpCD4XdfZXPRMBz2fRxy/2uDsWp8QmTBIJrael3PSq6Loa
G8DMycyQwLCnJDGIm7dvemjqJF8/RAI3XByuhzIUVr4qRFpRh6qlrvUszVLJHZqW
eWNGx2EysYpKC9+DoWXopl5l7SyxBYcBDQpcGMDbcTxy0hDnmmGUVBdCDb44ZeDz
BwojRXgc9+iE+q7MmgPIt97bO9vBfG/c5ZTDVtN6PDoJNaksi4i3AIYfcViY/xzs
LZ5iPUZgC7vBgAQ8vfMPrFdCTSe8CxJbXMnS+MG3VfOuyDE+ybp2tbL+M+oeO39M
q3s95ieTID8fs5FqCGbSnDsoDSQkA6K8QKqGY3SoTfmCFL6AyTKA9OgwhktH/dKk
R0v8wTE691cQHQOdPScfAvzjbiGQl0uaaHLN9vVo/ngED+Hr85AlB2dYIQ27Of8q
Nm+FQ9XSC5gr5Q1Ng7sP0iH88ZF28EPkgsiTcNHldoVkIcfBE5NJOCtWYSqC1lzZ
5xk0GkPwlY1t+c1n79oRQZsXieILX9C0R9TkCevO0Xk3Z5LGd6MRAG3D2c9xIQBa
yc+SUbwxgApVLbmw5vjMQa+/Rs+kZ8HftWdUHHY9zl0RrGLZZyIxZx5rfLsAD+ZK
ghkikFLrm5sT/kWU0ap0Y8NEho6ZA3YYGN5FlSjzPLyXR6F3UoNUY1XkZ3lfymEa
FxifgZj9bZb9zWO5oRlhBsS4RGN2JY16QreSbzwsa+86ibvK9qJKD0juP8eECMyo
+gF7HyvRtvDvjLxLaZh5K311wT8dK8NUnSVyhj5oPEEp/gL+DEB/itkC5AH+GkfY
E4xz4TMyfsnwMBrleJxdlhBfYAJryHLyr9Kp5KFTq2tFwLu0IrPJDie1NTfW2Pvl
66rvwa2M2tK8KAbdpXz/DJOxfcCdrb4yrpJ9ENaEN48UNETgUWft1mdt57jk30rl
McUZPA2fhwZP7YpuQcj57HMBX1LMvl0UERwDdVu3vCI9bjZNEFx5vZj9vgF8506E
FgAP8SMzw3YBzh2eW7MVTXzffoJOORuJ17yd8SyZkxMTLkQ9o3hoVWftHb5pJ0HT
RkwmY6bXahfwCmptMIuYMzv5AEAwtdfuM6rAJV54HmpWQMtDHlqZCX4eK4k1d30q
l6ADGXbQ5pfsAMZaAVbWonIDnBasSrh00N1cwjS8GApSoAxW4doXK8Mj7Yb7XZxj
ta2K7fhQA6twWcaa3Y0SwDnxvTECVi1RCgALFbrtiQ++ofpLVC7bjI7Wxt2dVZ3K
o7V/oWuvJuracO6/F9HsSX/QPJAOOQxoTnCkldtTHTDT6QEoR4Wpa4O206cw2fef
YaF5d4TfMtEwDX0PPmhhHfynEiau9FLLqq8EyFVWQwomLDr+I/jf5gbBMkVa/nYd
SW6Dfh3uLfh/Zp9UubuPSPN3/3HnBeAWzyagXZqsfSPw6fAp3EcLzCVvoMe8mw5G
EFmosOFieyk3SBWkjeJ2FexVj2uxF3+TT+1lE/nebOeyljerDrNVMWg1FFlMO4Qi
VhrDMGR9pfrMWA1+vMwvV0m4diu7GS2OfgmWvr8kZwryWMACiEnPF+mgY2mkAO8G
mm7i6LAKay31D3zErMiB4UT+iLL/KFE6RKvOkTlrTAssZ44FAIOOUYkJwe/MsaVR
TgDfJbxObdbE0VpgJ4kV+ptVLq84ASuILdkmIjr+sqloEDuOjD4oz0iyabm2j3/Z
syr4P2eNIsg6WUkLuK5ZTv8xJ9XyRYirKznmwQRNQwI=
`protect END_PROTECTED
