`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PcaSgrHfvBfYi9JTRyoKOOjBOWvt89ISyn/f0lRpqgM3zyFWKPFFeMrmsmov+an4
tupJWcNRhe0fU5PVJf3PCxsKxiIW06ypvEbFknImZ0+xY+TMXCtDT1bmv5NluATe
bGFeJ61ghM4QUmFyGwmrkSyH9iv8+/NWTaz+mNeJ03/lFRlUjRKfG880smpFL7jP
/FiNxxDYPGLedreNepLqoC04+7ClcPLbECbYuCzlu6mHb1gUGW3Zl8vT2IA8swkH
D2Lw1jAw3+2F66W8od01XtTRqHKuQEZj25KgPSF56ukN1YNj+ihdTVEMr2JuDJgr
n0A2m+TgU/GEj/H+9+VFpI/gPzauKoOB59y2AljQWu4RN0RX7zIjBpVI6S0qVQhX
AhE5nZEU2ACJ5oqSgUTA56uSuX3jsAENzHTDMdwCMtKoIW7wl6cI3Ir0BFkZl1Qe
KfdusBmX4adhHpv/VJN+rNnGIcE+QF4z5626bea3McIxjIMn5OJ5PYnNWz8dYubd
4FvcA3bnacewRcSvdvzr1bN0/RsQE6uDhnwsqKdnaYkzyNez0Dk4r7yicR/VVTV/
DNaeG35SgtWdwA7aGHC0FmYhR3+sPkOTM/68troOA3XDNtmOFFm6nbOzPUoM746Y
m5UDZ/2pJlenuZ9sSkLsow==
`protect END_PROTECTED
