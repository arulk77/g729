`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGHXgYtkkeCofJNNw/HngAZW6Ovey1h+iHa6y44FmAc+
jLMO3a6Mw8uNEab5Xc0HBJwGd6BOErvllJDYdq98pNnwPagX1d4taqMnM8ejRDSk
Pmirm6PMV21rZm8eGHfZFg+X1MccJxukihJyIOcEr4XhK1ZRj65UT7GfaKsFpIoM
/B0pUAO5ngyQcdVZ6sbLEvjyaxeevgn3DH49LuIwEDwexBbxUxQ9snHyXwLeSXDM
8Wd2m/7jOSLTmDOCMo8URw1XXeKJ+DV4fcyHTVu31M5+O86MasiyCHE7mL9U9WBF
EvO/g+1xKIuWsePoVhrOZSfOeVf3qiO9BfN/GhYWSiU=
`protect END_PROTECTED
