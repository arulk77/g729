`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIewxqIZaTjjLFp6G1YWqYY9T61Smkm/0MDEq1CeZuqz
j8GPiCnRp+6iGHNylPtJDIuL2ISD5EA9vSG6/bfYYfg1Z49DF/gqVQbA6EcRu6Rq
MD5oZkycoJ6KbvnFZW/0XhPbKxBgaC35+lEWzQGKWuhM6ln3yZPdr7kNK8g3Lz3W
FatWqa173gHw+K7CXlEmfgr4zvJZ3kzV7yDFJBBxk/iLdox277kG4z1AldHc6Au3
YIJk7YTPLcERsVZ3LhPWAm1YttNNdhfeUwOZ/xPXTfUZ5apJfG9KuMqC3nfulNz3
WTeMx9HVaR1U6KWsyl2fea+pDT40HQU56B3mXC71LdA/QZouSA0ONpdTlxLCw5WV
pRfuGPuuICpvsMyalxoyZ8XTfYA7VR9qLrSMHKuQlRLIEd+Ei0qf7OzG6rjQzDdt
cJBOAqQsfrXlBCnklHGXIPhKrv8id+yTWKwO6KGNl5yyW3w+RD31HY8HIzVoblTq
EnEXDfF8FKrQNDyR/6ThsA==
`protect END_PROTECTED
