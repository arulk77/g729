`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNmWA2S4Yt6vb8LdI6XRQ/eXzoaoHEOm46IEMx7ZGKgM
Ocabf5ZyRlNuFvNvzLdjYLe6X3zuZNQsDuE1dFNXAnNAKN71EWVn3W/gk6YHpvJM
sWBhpKdkG8p29mCNojDEItJCwSCuFZYX/E9t5YDzeEGKxdl1pTMzXGnuvtIVuZMO
M7djRl+D4dlv6i2omanXPbQS6peZBfSRTfjYIBVvl5/Lj98j8nBQJIqK+6TbNbs6
WrV6lOJJsA4gcJqQSFXq+SDmCAOrEaQQIyuzZLunBJGM62YESWaZ0zkqCmlFENnf
FDIb3vtWt++6jJM9cILq9R2ff3wtDzhOptUS2ujfuTaL3mXAVE1hWehhZWVcwYJH
`protect END_PROTECTED
