`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDeX/wnFyHVE4sBcNYBKzlsYPwP+Juje7dUDVoeKJMwf
24TRo0ZZN0ZYcBkcz0bDARIkoK3xfN+0E3yCeIcPzCb+M5l+kxn9QVljJuNJf+C5
wNGL4dgINbqGyG/m9qhhWu2TZPJirUqxk5El3/gT9PREQaF/ZL7x/8jsQ+XfLriJ
yIjMhi9n6uYfcwssvPqCieq1t195YRZoghZesNUSGDDPMYZD4Np8ry3WKvaTAWq+
JwjwXCRsChOaEBE/RmMXoA==
`protect END_PROTECTED
