`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
v6DFwlVhfRJAxLw2wbPVwW44wmkD0YBNbwsjwsxuBNRWffFSZBj3RuOx3k5elKcX
yWbCARtjLu61oYFxii3/rbMVlQE2vCp7F8r66/E8IRsxKHck8euehi+DHlbUQ8MN
ytZYSeKvD9XzJhej0Yqym4SLglP7sgNdkrwxqN16qRGs+FBWCCg1yXbzr3WSE370
FaC6RNqlwBbm7XrXnPXxDwKpm2VKPpw1T0BKnSd5QQeJ6KSSqBMx6p38sN6LgDc7
n7Uj1C6gPsbtHiBFbCEtUWSw1MoV6wlVtmoj/ZsGYE0=
`protect END_PROTECTED
