`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMObtWgmy/AYDkk6TJ8xHpWXvfcyVPIb8aLSZJTenDNl
hwDRGvP9w24FDEstLyg6G1cBENTot5Wbx5bZ5mtjR1FiaLyTYQKmJxYs/SG5eUig
fsyPTUMVe0WW/iPpnq8/MeZfxLwTLGP4wbOXWBtjcp33vB+2dI5QpzNJlSU4AmxV
vHiyN6d/x+8IOSvgKN9KoVriBxs9cmv1zRm1AelfK6cOtJUvQt5tliKVE+lTO0g8
D2V5Ahtndi5k+hKxlxaeBA==
`protect END_PROTECTED
