`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBP+Dyfj254qk/GdUOGHvVV0efaHGGLhuil6EjN5G5DH
8lfVoFrnjJfBhv0fAvNQ2jguE3b87G/upnvRpiXrZN1imMrBKgEJvpkkL1JQQc+A
Ng5pcn0z3Cu1jr09Pawi2SNVoUFhvruk+43tTpL/Pe0SyvRaRdo1j72lLBFSpZd1
04n8JNiI8TEImHGWfoil+6NVV6KojbKmoOpDeH3qpWrWnTXnFT/0q5DJDe8w/mQP
3d5uuKhAHUBQCCgIR7DnU9PZ0DrwnRPs3+wGtQysBhobt0osZHVaFsnPUilbe82X
xuM7solYTqU2Mv1W+ILPOGgOZfHkzdQoFTwZUzScVwPq45aziRg15pwUrPejResj
Tc+zMvGLh4AYETn/ld/lLAqPcSh5pBg4Mh+9WaLqBjJcsqd/2myDlhWgb5fkBmCm
m3TroQRgruDbK6IgbbHz2BDTsFBBGalfV+gG5N4rqmWETWl9hUkhvgGVJ8RgW5V5
`protect END_PROTECTED
