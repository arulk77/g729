`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveApucFMuzKRDVoNYNVevzuxYjpzOTckxZX3WGVLtWCQf
HRSZU0PX7eqExCWFZjtufkAQZEpy+kjAxnIfKPNVKc5KBtUQcWU25pqHt/jih/hR
x9WCZVnNyeVvO5TrLGqRnHC2dL9MYmSccArT2QDh0RUoJqCB+s+GSRo6ITe7C+yb
aJO/IYDHaENUtNJ9S14fyjcZUFVUDv/0f9B6RIPqFwo562SVBxD9ouaGJTDfk6H1
bve+3j26BOEe3fQps0zjLYRSVdiAmtoo1jaEmo2PxPyrhupxAgnjTvNuiVipcw25
cJK/artk//sbmYdW/h4nQ68BAbpNn16HgfIxxW2myaYd3YJKyhwtB3NnWY6uOVzn
5j+nscJpOOeotlD2w7QfrrAhkoMTAuNQz84EvBCXw0/xu0DOpTvxej5NjR0vx+JH
9+imqxCBTaGLRhGWjpZfb4R2UzwER+kvBvlgUMan+sIDBQW/LfYNZ0bIsF7ZjuRb
PBW2PMySU9KRuc36yxHiBbXrvRwmTk7BmkLi1KWTsPDP7MlWw9KxZOn1ReyMpDW8
kJhJ28fJXk3On4BMgQWza3ESsUuP1Z5QHO92dixwkKwMv+dEdeYhF7cuSVYBwYUq
ntQIA9+IQkXjMuB9clYAt5B7ziUu0oESeWBhVqnL8aCvWLpYNek/fn0oTGhEA9+3
OqByhAmoTiUnfM3gHXFoRfjMGDDMD7mex0KePJJOTrb6el1xo5Jl2hx6EWSF89re
OFT8/hRqnXlzcnmeVRQSsAALy4VAgCySDzY7RdwUL1maryICE+wrMaCjz9G7bB/z
VqGQmyLM5gtbRlPpYNPjIQdk3J2KN2dgw9LSO+riKBeUgqomVQ1Lsq20qGSCx2uk
qND2hHzM69jOUZVOoYHUwaEKbvAodsFw1rPJLGT1xTJ0STz/V9iAi0wKz2H2ahX0
aw1i4Znmh+5QzMkrNkZz/GkZAROIeCBU1B/CZnK0j8htZaljuQSgTH9QQxaJJw7i
l11JMgLUEiuTSne7c8rVgt1RhnxiAerMPGNyrlm/Cw9DdIJim2V0E83SLh6VyLqs
Ik/hsklsPgj5Xh8VRvci4i/ZJT+Iez3lvhrLcAp+1Z+RTPbZ6F4gE76q4eq2wsFb
4L558ISkLN5Yrt/2711cV41d8rkPoiXBvpo6LqvEn35ssn+Dm8g0Ydsf1AtgifwB
7l3F8ykpTfAa2k51zDdUlabCPJs3a6rlyWe28OrNeSQl0w3Krp+4XOM1ssVlk8UJ
53N5MZ3Q5CscWiQ+eeLzPGA1SmtWz5H9GohQ70EnqCl4NZaJS8Lmll7m1e4UN9zf
AIfDuxwmGjASjYSMxqH6+abri6bebJkQodNNwJOCbCJ21Q+FRpJL3t7IVZaymXF8
EAsXi1fAJD7ZJwwePiohq2rntx6MK6lbGc2EM5JWsEakqUPXB5IdpbvK5G6NTeov
l1NGdfThmZ9/B52Nink1EbC5rhQwfRnWpZqXRj1xjp41thVujmNudW87hToUSHBj
d6HstSBzwjAol1vIkd+c09wcinSIsWjLkwpLPDB3LbaOPlY+upmYyJYJhjLI384b
C0Xzxlh/BoBEYp1SVjQSdbBQoqUwONfetblHa+7OkINggcF7i4ZMxSFGG4Nulb9U
3BR8aKScbMrcbjEz9zLl++iwI+S8jTn+en0iRXq5s6cAMuv/jtTgebpLTS/G/1SF
4y8jdgEWmKz+T58n4FsS5U7DXpYdd9lMxGHx9TP1ZVACVCndGHvl+6zPbNmR3M4h
zXH5Ggm9+dTjslKN+lfI9XuXq9OpCtS4mV0GVOkZxwH3stG75OjYeQrWJqxCfUhU
Pxi298eNWO0OtU34O7cvD2mHIku1I9R4k6nTgssLGNkZzhZA5ZfV1WQE6Rb/0o7g
qYgtPvgmxjZVpD+oZvv8E9iqD+9UtByv5BkZBAVhdTbBLsiFwHTqeT3lgPUmEZAI
UUPjQ/w2Yu2+dGr9rHCipuaG2BBVgj/oIkTbLehfHYwdvgn5Hz/QQe9HgT+4fAQP
8z0+RW1q2NcE7ORs4Wckh2QgRlQ6lFx4uQSsr4Wk6ERr4KghkSlTmaXjXICTEu6B
l4nucVWyh2AAesdXIAaliyEH9/0TsikOV+pbvbcWld51FV0PsAwxj/q74RAOFsh4
TOA1H97Z2QDl2VYWAbBRLHN2MlGmGeDMwHQwbVODDuKv+8H2tbAHwWHKmO1qG7DW
ptLhDJZjcYkGUj0sQ+LCc2WJu+JfKCX3cQJzsWGLVTtmQkqnwf71TGSNkjFqg+sp
t8bEdL8iq9zXF7o/KW0bK3iNncPiaigqsfKai+Up+QqzfYdljclx6tARdQCuk8Nr
FwEgGDR0/RZ9y+EjmigzAClXAx3ljm0xUWNcdgtsrH57dU5QXbZW7AbOkpsVv7mu
xOyFNHVWK37GcWjxymzkZRphoGJ0QikzsxcUfXzbzsT0DLJsChJR8hScblatkPJ1
1Z5OsJi3VIfxSxdyeKVNigiI4u+Gwd89TNzg2GmsjemZERH+XxpQpX71lGNnlrsU
5d+Y2qQ8JUljBKkDPapuKrKFPZKDNy1rK52DdxFt9267Yvb3nI9Z5Yu6+7LfTlGS
7fG03RuxYidl1wNq5mb7OmkEMc+HJTYgJIe5G++ojUQeQOm5+/6UJ7Mo4QWdVgSx
1796NXvO7O019sbxksoX60iviFAa+4XT+x9wS5nug1G5BJu7hfWM/4BVa6nLXu6n
tOPtyKMJ81ZP/NqUGsaZarioDnmAffTgtGOQSvsnyHXExA1Iy0/ZrTBQt6Qg8Y97
j4pGcCBHFjFQXWG12ehEyNFQ4WFEB7PfBA+2eCBA5uAF++D/PBfLXLaoUyjj/4O9
9yXgcJIj5l3BoB6jqv1NHbrnhTNRSmq0ijZf5KIU4GSyZhmHyoqYpkYVvIXycwtt
D/KjzgBeKLsDOBFkFnNbimh/t2cJifIBSMGZkQZnhLjLRjouAXVaUa31NsG1So7p
ZDnXMO8zpp6dh83x5Q9JA/qf4P1//7AgHuvl988o2miwmqR+SDtwShMbfXmREqS1
V3Flku/cv8L3MWGdjGfiBaNL7QKSsrNg5njAkR+XlA+H+xLHPWfqHzWMoPeSjxOJ
e8Xbw7aWusD199UgQbdIxSgV0kGDJWhV1yciUoZBS5j60vQaVfxg54pw94bY51cD
RAYUH+dByp9n3v2yShvuROyUQcsLQxnlTpPsGPozKUERHge7t6fuVemAXPiZS3Ik
A2SWnGujgfhQ02REeOqosoInBpY1+0TALQTsIXWdXBfZgwmqr403gSvr+mw/alxu
1gCmi7g+Y2OYmo1w6HC9Soc3DptscARRxIkebRl3noxDnd1p+BX4BN9Al+TE/2pn
buEsOA/lCxnxWa8Ycj/CZIAa2Sq8QfUTKUFnKyFTL9LqfpwiSZqnewbCtbebArpq
SOR9WztGvxRaRbKS7jcYn9o37/IBVkGnEOsVYQM5C9516F+CIubPIeGDf/TcRh90
CuKXrgMUseyNU1VSYFlFanz6w5a7Np1ZxLh7Rwqrxqe1/VJz2CzbW61Xx7lmd9y1
Wlyomw/AFXSduh5Wmn3VVOM7iZ+G6FKf7jcZbGiuD8Wtk7x7ifEaWbr3bjYlf8we
ytycY+2SASPPduNFxWxPMiDSSs2wzCQb3qomlEp5lf8HUXietCAnAkyKXtdVHv/L
RugoIMz3W6pZYLIQ0r/xHYc6hBYiFHwRO4SYrQaAN2k9FsgG4Mw2vWRytwvac+v3
uuzicHLkxTLouJEKhxGzl62Q1VbwHFX2tW+omw8lNeDzx3snQgDmWje2wGRZ3Zow
izQoytnlwsgLrADG8WauMB/liJsfnEgqxmCRX33fjkyYcnUiqCnXuevGac+vuRe2
7jOCHJwtUtHpNF/O1vhVP1cS+b5QmL1sVf8yT+m4YFQP9s+Qxz8EgTIr1E9PJ7KV
PJhKemP3aSlqYlneWXE6yYlBPXcsVkTi1Gc+gy3FU453IZ8cYKD/Nkrhn+ezK4dh
0FtShBRwTZA6TrVglqeQefHG18VqXlsImQ/Q/XuSoMr4w934RisnbBhahIIst/es
CGgkcGXbCGzgcA/14Ov0NRkGG9qTZeIjWgZClazV/rWhrpfmkx+DW/sHNrGrUoqO
G+r41vPDYYotCxrJtEEqg7MtbCDNacGXBoZWs8opP8lFnCYYvhjUTA+yeElDyqUJ
bodj3DTPYQJHvP8mx2Ef4KFClfhGHqtzz43txat5wCI5W10SqHVpsmbABklGwXWM
a0KG7oMw6bioIxn1/G7/IT77a2e8yrfjgulY8aVdkBJScItPHsxUZuGO3KSmYTKx
J4YgqA61qkoGrftqbBNa96ogFUEH3VMEqoaIDUAhQkVBu/wd/debOZidB555UXFf
heFIF5wNr6RzxGWVrYy9SezHoRLg3w2VIPzT/m/5bPLG8Pwl+5Whd1x5o5KpGyKV
fWylgwZG7OtiXNazTXCcx6u0YXiqRboWNK8B5tgKMfOjYVI8hnH6Yps197T8mC/s
YwZcpUIucuycPZUkwyEjdo8oAudImznix/+oaAr56zmXlm7M4cWdOTXnCmyyTMi/
G1dH/ZSWy2x5/6S/DOmm7XpVO1Da7aMxiRjGylWQxy30djX4N+sjtXmLG6Q4/niL
xhpNmT7AhPWnN6hcJWbFpXM6JmYLPg87U9qvWapr78u3N5/QhQkvpfFyg3bgahJn
pZh0NiTzL/kW5SBAlf6RZk5W9Ni2yGyZIv0rr8lvdrfzvq3HBCIl56PlfkPzMXTo
kTlicQ2vo3MsHXNBjmRG/bYh7TW31vFSRRGcZ1atPvWFpdx2aEg9q/UCegYsw1fD
ZL/LVZW/6BuBSHnr+zZZyvwkmBHeuVfy3ah2SxaOqg51no+uhMS9pT0D8pViPvv3
AbJ1YTI6CA2SgXq1s07CYJ7qKcpMetGc9HVt0QWb5N3MKhaLQ0txc+uQxoymfOlS
xrDfXhv2J0V/Sir1octie9mBaHTFxjhE9WTP+zxeLsL1bkI0npul6gom56sQItUn
enKq8u1BKtdkom4b5KHi56ivwWY8BBD+XTAAZibVJaPkE/swZYVMqQ4UayWZwdWl
a9Bpe8AJSGG5jp4ZUgosidjUtn1D7deOF1gPH8PHLowm39mjQRL4LDRi4xpu6Qq5
H5S3hUmUDkjfLdmACKTf8gJMJ26eTbqRT1/cO9Ya7SaePV+a9nNjoMdl04EI/atW
NT22p0mh16nPzEKqm7MXJG1oN3Rry+R/G8JFWfvxDfbr+DnBWOih75gQrC0ZhBbV
5Y1foLB9M4WNtMlVbt7Hpmu7IGJKsxo36Tnr24e69lwv2DD8mn4YkupfbvSSZTYQ
7OJxAd2LnnPpT7v339vVV9F4IL6aAkpMPVoB6uN5xx8ogG/6V8CAMREh6xH6TbuL
Yp7a4M6OGK0UVcG1mYBi72yTD5iLrYli8cl229DIYEohVkyQHSyd4bl3gTw8ZJQ1
fEAEIYWnSLMQt1N2p1hXo7Kg2Jr8hH7VShq2F443og0N59qCnqB6pKvZFpvPC99O
NDSgw9DcZXNZQH4eadcb2t8m4c7BhCzJhtwahkpegl3scWqGyFLqGxId6Rbrpq5I
t1RXdUfyAW8EsWznvbQFkh0xi2qG+F6U5HkdKvxp3KdlP54C5MmyaAlyKVJEIpVQ
UsOHGe+CNb3SP8nLFXN4Bf8214fDjEWsHzoI455I2mpofkwXwiT47isDffQ2ZOAu
5zUOJidpOvkvOmR2NnavTYTbBnG1ZHqD0eZmFyvB19Xg7h8g4i+FUWdeerk7nU3u
/8oudF0GAeqcFzfF4WNeFIC8kp6FIsoRLOsEgecZM3wvTUIjPPd1ST5hrTsMOLG7
ynnY5AZv1deM3nKgVI3GGN5HWy8iMRvYIWbxYohL8fVFliMat4wtX6uaECK2p79v
DwaQucBi5ukDaWF688JYE7ssPB3BnuzlTUllHAJjYUCsxqOButBC0hkzI3kKNdfv
gfMdcqnKOKa/Mx8VFmyE9exq7ioezq+Y66OXyC+CwNXOxVnHMSKJJDgB0mphoks2
cwT7q1vNJ+XOH6XbB/CbYmstZ1EEY2a/3weJlR1z5yMSasLkFClF1k192F1qaVgU
tPUS990grY8Yfr9/DA874cqAs/dEVwX8xKe6tdh1g255ee5ZLcdbro8S0uA1WaKv
068BcHnh0WlZTnv/AsIMqvNQPNFxk+t0hCpeaEOvNUYvR1r83icYxnHMnqVVKNS0
ug/XOBWBIlsrLlnOMqro1fyu5n0QPlR2ZH/Ryg4EGutA7BF5rwRP+36GIaUcQ2sf
cZjkfnGYfhspq7jUSULEQI/7FAHDZtuxgIwtqL93EPvv7ImhT32zjqoFOH0M5ul6
Pi0K52KGuIl+DSC8RIwMyaAk27CBzJVCpPMQ2PB6QGtH4a/qFHvMunG1g1uJbBwK
VeGpnP4dG5GuLtt1eirj+AWOFJ5go/BIRxi5d1erYmnXWSWQ3TrKnpwzy19AvDiB
MtoKAr3eSeJqR17tAiulmXDYUGNOrVodIKEkh89G0utH3reQ3yw0igVFHzVGZKKt
fmczsr5c+hsqtd3hTxqMqG8I3saPIhYWivqvRPcfUqa+AvEcu1p5acdPif+LGfs3
K1ik9I+u3qLsP/c67+J+SJj8S/ES6x6qwIrvZIoU0isFG/+IoC+uwOwZftFO5aCP
QHxtBHsz2MQSu25zbIUdkhKz5D8olFYVKA7/OkBkkKjc489HWTkCN6/nbG0iWjZV
bCgwDXg1awqDDKOho0oQSkrg8ywiluXuTAmEdG6VaNzDfgk7OSe1W4nT/tcneh6c
07t7NFrazbnUFOncx0tDDW52gC92gr6QJy8oWhouweiTzQ/tpbcdyo75y3WQsw8L
nAaoVsoIgOs6w8z/j9jVKswIhf3YJRLyJ3olivT2oCvzZbjEKrIwBV7kV35uXOZ+
xS8QeKftJGwpKiBwLO5hNEJ4qvnGOoNXavqWPJFTbtPRG3+g/QnnFB1qnjkcFL+x
TjLVAYUfxRFemyU3PwEptV+mPo0qED6FoxCuhh9DwqVxROsN2iox8tGjB7jt4g+y
JN7pcrgan5/XoMyRLj/78ccAnQGki2Vh0MAVsfAaXSouZCFu3hYiYi+o05Q20QEX
hvPyWOd/9SQ7vfxfccVsQjIWMETm1XMdPR78if8iXzSXa4FlfVnAEx+ZnJTcFogH
9JJnURPTzL/7fF2PPMQvA2brMMKaFU8G3vCuHEquik67AhXyOEmA8raiIDal4tRF
wtSQsJ9c+yUrqKqR09x0JKO57O7G1nGBnjf0ByBP+j2t+9vbsj3dS/Tl+KSbpzjJ
BPfEnN6EzEkHUtbaT58wPRCTNlwAmHuup87GaA7nEGxk0uNoKqeyP6m2UJ/HhWRo
/VsUsVwWlW9vLidnazK6Ju9JY5SpbGymmasrw6IJn5AkB9XsoTl0G2d8yuhas2pY
97d3ef4NZrX/M8b0L6ym+B/BHYltbP5dIwNrG3Wk1Yso4dpz34kcAdxroLZJB+Q5
raPChozKEr7p6BOdoSDzg7Yrd87eD6y/htG+M/TRdacj44c6PWY7fLShtc9goWab
8SAXJE9oAouTC/1Q4VXlhRNSQc3/ozpJrBfHTFpb3qGS9k+4nPNARIaJnkYp5vnK
yZIcQ2Fg8HQAat1oe8uh02XwenFbpIreLFsS2PFK331aIunfDU+9UQtFmPP4Ojeu
NrGP1RI4mbRMSvQs5129UFlVNWvYbhzsJ+pgz7To56CNOGUMp8Dnpn7ifk1CS12u
KprFrLuO3Elg5Ps6+hThOwkRSLupuqCDaoUzJxAVI5LCNi+u1GgtiSrKhRcGxdr0
iMbBH72TvGhyUyrZCed4RX/iLDypj5zK7VqPb1p4zlMUzYkkcFXomJXQQkCtisJY
ed94RI55DIK8eYYUGnm4VcfvK5LYzvOmgOp2uqIxcJHbaby4pS4Q2+sGDnLMIB7M
w0E7bxiJhDYxnEFy1gcSWRHY7v94yWIC9Hu0SjYn3Srm/RSgWXAZymAeAkAu/g8E
dxS8uSZwMsO+UucbiqFBfW94vouSiE03bDwjUXHfDG71K4HapoHyco13s0mz0rny
xdybeI/ZKJv0KzdpTf0JH+m389//Mk0aXIP1qncw+Cz6nkzFqNahjlftffqLAodV
8M3dry4QuT629B05UE7RkgfwrK+Kf3cZkDqQJW0Ws0Ht9J/X6yZT2TI89/VmoVMO
NpiJqSzKrEykgUrA77o2YI7hCoWLVbDv4PqAGhp39GNgC0YiQuohnpzm0SPL21nF
72Wi2gukAvvdMViCD8Q4yi3cZvbmy7uzKB9VTrLGHCCQT5gK8iubkfSbKv8dV1o2
5Ry+Xz2P6mhqNs5PQ1zFcvY6p5eGvIBuqGJkJf+Wl06eFxdus5lTu3k4UuaHSnr2
H4EHEZraBrytfMgWIOpGOk1DUyTC23qFgGDJ0EC7zKo6rVIiON+WKhcyrjQ/jskQ
a5rxbK6pdo8BPBjv9e6A0INIBOA6tFPuwSwqyFacNQ2dj1HQwuNH52jT7JcFVZ7Q
WzRh575ioDWjQ25ttQ+OF/JZFwbZCmUKI9mtiCxMuY0+CnZsyd+e6yleqZs1qfST
xTRW8J+5r4VpivEhwaKC8D1O/0qp9y3AHgrUaPHUZzJxKMbdhaj4jqN2lW53xCwN
VsyZ80JyvDHetB0+UphRpK+fs3WbEKkAnDOpnCcZCcxjC0rTM88IS45TC6z6nd7d
Xvv+7USSRq/TXeEFDbO51PhR0gcBIHKp118Rz/S0hrRR80VAkjbdM7XvEApBwuwd
2dt1MudraduUTGMzoNaMwS5DCxmAtyfRB2Lc2QoFIrg/0FR7h/ty9c4dXrDQ3G8p
PGeuvQJ8UaSXwfCrKNAfMezBSasQV7oQNQW7jLBfkwCO8oi94FCLs4qZDPK4Hxlg
0KoPbUVLr5iC67gy8C7s/106S6/4i6DQvsCTWXmZi52HEGhZlNR68uuYhFC9WlUa
Ha+bLk0woiVBAXCdICV056lvkFloXD6nrJP2WrnuPErBxXzk/GI0w4mm1PIQX/si
XhHTfTbEOHQB/baFOyJrmEvoi/OOL4jBwVNaIfJIYnegxMkSHBLsocwPGDNYcoJC
5IwZRFPRVa+/2tjjHBXs3JTGRExaNFfHHj55tkd6kZ2YtuN4+vQrmd3+gLwGS8k2
CkMbSr9N3TUWv4MgjP23GTze8D5t9197XPmEEyT2jNhFUv+Tnd7RCmWD35RXxQs3
eclczetP5NU5qaD0fkCuOczKKKnF1LTJOI8GpbSJadHAMDrJ/+O1lawff/Ahv1qE
g9uOXDN72i2ifcK3O7f4YqQe8TOl70O7BTR8nDojthMLLM6vxmIUkOQNFjS5e3tB
giaEQvq4tGeMkf0aJ8nQTEq5nVH/mtbstdLEuddTB88yiCN6+4L8mginl/eoYmaV
nTGVCKIL3CCE/tBBx0qiuzAAhYyo8657rDapRVCUQ9nRgyE7WZM6858Ki0WL2TAP
gXzd8Xaq2exHYLIob88iP658gkjeACfqcH0vXxhFWLWu8/b7i17JcKPpgnRbo/0t
mtAjazMXR9e5JD8FF+QpG0b2/WVtxhOokIIgGJkKxXc49aiJjG+dIzlpYunLLFnL
9SP5gjzrtdPni//zCC/8LDtrITkfDX5ZbxUodyTrQr55PrR3qByWp2d1BER9v6/n
HEc/nVqTxC3+oClag6IM/+Seq5k5uOfTY4edcQbJzbk38e4jSTEDt7UWt+RSmgh6
tx7phWcwQcNEtI7g4BGIhveEkbDMAVXb+ntaRF+4sKFFYFvOC/ovf02ZLnolzuTd
gqF7p4FnNB1UNwmozx9KUY6077+ijK2FuHDHvJwORGHGDF4Lo4bbWHzN65gW6Zhg
uxhzhJRNSDbG1ZLhVKSSYbggorjrCQvauIo9UvDyxtvoyuIEU+QNj3XF1YcKdg90
GdewNfe6CxrO4sz15H2G5FG9LUbeKBdoq78c9HhQ7J+KTIHb/9tbf53qWkX8E8qu
+mUbhVYRP61z87UsTSKSNaAyEwYQgMrid65h3DkeLKydW+n+8bZiz96hchvpb0Jc
rDvV6BfcXa5SQDwrgOT7FW0kTqXz3WkFwX4dl7GXmRxC3LlbE5l+9iGYD8h2CS5e
ausutOXLUjxh1oU8BYRVX78zs4etoZEeXCFwhXJPXrSUV5F8TvThIPUs3Cmn2fXy
2LsuujVV1Imyl6bZsshkoJDHx4o+CF5xODeOrpjpkjyJIKijvYDf6bjDV/F9m6Xt
kROhjVeglhx5xlIcfmyGdv6DVWPZkEdnoj9AaglXpCVIx0aH0ZVdNYBogOlspRIq
6WKZiiuCh3E1za/XRcWa6AJ5Nd6Q77PhNy1DHCXi9466JtQlkJn3Y36rnykbXr8N
8+0OH0E9GYSX0XPNX8cKn9aliUEZj3FK4idtaim4ERtTPTuCVHtuMelNaFIobVil
3nk0CP7oPrI6s2qH3TpPptirqfd8vl8AsyHdvcQZG+kPSu+0rXbDR1sR4NnGmYbL
/hVzIk4hbUGfsxkiX+d4XC/jRMZz96whBTm5MJNoRGpNVC5a4MoBDDOS2FeTpDmj
x1sgEg/b6G/AcBliMUBD0zBc9a0MsJII08h1atSlaDuJxlMWsxHTLj0+0VMJkqJd
RVTPIOGD0cIsw0EgvIsssnUCYTcJK+fDG4wCoXgDjbJ1uX1WefMhQcJmtIZGGi7u
wtJcgfrKRn2fGO6YqVHUwixe4VPJf0Pt0RMXTNI2koWuJfgJdK+32At3t/1TINlS
hCr/YmGXD4IhaGG7iLXG3nEdQuOneMnnH7FHuwd8y4iLUoF30EGa8g9aHFspwWfH
zA4dXNf+e3wdCnXf3CztZpkUy73GaklUSyyyx5KY99dOh9zCGu0mukEokqtRLnWn
cURugXIcRrP59/5o+WWF4z9secoMzkJ8797OEe5UME6psj+Z32q2kDs9lkOYpouF
sWoBZOFqgh2f2egk/zqX4KK5IfRy5JzL7LKQLFG2iU/gXlfEG3btUCXRZ5MXike9
TvLjoSFE9yvm19TTsBf9xMtHVEhScv+cF2YUix/IsAGDvoCd6fV8MQFVT/uTYMUB
wzYUJKdJ6h3nqPJSpAm1nsETYsZ7E8f+xrO3hGxAX7Uq9lNhCSPxVRnoffeK0mQH
Ip6TTtegCCEnfiTb2RozSVAperwOwPfpfdZFxF8iba+2wh27p1mT8ZazwZHeXM7u
gWSIZBK1SIvuZ5Ic2NSkP0DcYU4aRNYYZfPiHU/mxZhDTr6M4RvVv7J8yC4yRhNT
E6sm5wraqxd8/ma6kD+F6BJah6ltojcRakJtBh3jYPiSqow7aUAA2AcX1yoadX6Q
yjPeVf4IyJLXjBizgB34V0lijjwLCk1w6BBaArcjX0PmPBV5dxNkvMmeGl0eW3f2
VFBuiK+7PyoOM3C58IabRrl26PKAEjD0Fp6+vrMRybV+VcirmnCYYTZg+7oloHpu
pmGalzOhQY/AVaKbHlE/V6lyBMwUlLIEc0NNMN3LQoLj6AVdmNnPRXZLvkKdJ/pZ
bj7MNGO1lmr3Jfbh97MyA41+VPJ//nVSfpCb23p7H+FSBiF14+4qt9aYHzyZYx4t
20CiwEtPCZ6d06ASWAMZIRNFsaaIDvn/+pzADUajVQv+ekbczMoqbl2NN8hv522e
eL+FhMc/i/yHKO4Tw22V1OsZIGH+agD+TxHhV3TUIoaQzEIZ5sWmXqwNVzqeJ++e
IV/r/NxL2vIeekPyDZGZAoV/F6H3EmryrvDN1YsDmsKZ6G1TLe70h2FyZamWSPP4
CbiKnqi8ibW7sxq5bqaNmZvzjgm6E/sGc1Eunbqcllx9+zzchb7CGem/1yTLhlh5
C6EMS0l3BU8roxg9RkhrrA1DGmbNnRbG8NtlCitt4qygOCqKh8ORgH7MHHOvoa3I
8m+sgWghC40WldtB8XVIo4hdSvwW1XejjsyoR+SILSAh2hs9amyuy6M2KDIcJQhE
urFMShSllnanGCg6coLalmwT+Jx+t9yQXA2ThyflUSzP0SVHXnIwetVLQ534n7ZA
H8QZgZjAyDghPNzbNaQABolJyEmpjhOHKJ+4b6rZnZAbRosLh+5BDB5xKlHwEgWT
7MvT3yPC5P2Fq7UksGKVUo+sa6wl1m/kaG1xR7P+siWz/aDl2kmdFh+4adq+tAEk
p3/Eqz/7vk3k9Mox6NzNPZEE6r6KS7QLRX5yLykIMPudUr91x3n7xlFwjsBkEf9J
TOcg9ZWGVfUbv4DXMRBprJnxmW29rbSbbFALgBB+wORFOgavVCY5by9peo+m7blP
BrLCYoF9k6Xq5JTho8690XsyJw+S+pvinUo4hXTueL80YQev8hWFko2mcHl3m4ZE
wiyrmAS1NF6oFWtun89Mfuu7lOKoyHhUMqBTaOcWZNCkZnqeSEhYVwg62yFMRJMZ
HLrQAOpz/414bXQQ4GOab1TIvwCQCN/Y840WzG6J9TQZuAQpLaiR3RIGt3vjkdw5
FSAcf+KALDlVZpw223hg0gr3Wm7TSGgEKoXR0MrB8sEjyv20PFcHlELMzr+6lWmT
+zOb0bAOegB90/x4IWAIZxmRWAIi0ANRiDcR6u+ewlaw1HdcGt5mUxbHp0F1yO0o
IpTlhUnk4m8v3jOjYbWGLex+ATP2bmczPpglWWVFKCykHdgBYET+kBBWJIGvMOFm
Y5hgY3pXaoohICCibIiSAGKQvqw6yi/03WfkvMs6X52OIURNCW4cf3cxTDcceARE
KVWoQCItG7TYzkMEncP5hVqHh2cYdIPBxiDC/H85qnXtQ+RklEREzLI8QdFw5Z7J
3FVUPlJtmVaKIG3e+7K3vk/T8DoVnjW6ZpXXJT4xcHxDV3tJoY6aqwgsAq5igCD8
SbvbFYQZla6UloV+7NbONZigUkSVrmoURw9DrFvq7TiPO3cyt5vFXBZ4kcYyRLoJ
PrAN2PmJw+opB5hYyySAfk6ywnE2erFc8SPtJ63YEsF1GhdDCH+Tg1lXdskVYag/
6aRR5mV+wmNH95wWvo0IIXKikx+1Kfy6Lv0f3K1qDNd47NY8kgFO5wIELzTNCrtk
08n0YILck9qHTHrhF6RDijFyz+okKaNqAKkzeeVzlN9aUHAUBhMWiEgy5oLL2Swl
K4RYIvwl7pkf8uIIjwxivNuZefA9WbAtPtKuSKvjC/lom7w9lTgdcT+XvCGUq0zE
UQ2KP8++3Vcwxe6tCmoqpw==
`protect END_PROTECTED
