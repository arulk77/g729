`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ky8uZEDW6lvmS8+b24L3FRFILHdrupeePeLZFF5jRpxC0anmDDw+7xNY2qllsSn/
OYHTK0305o3SCaKvu7Y7neUfxvU+eSENNjbMxXd+qnYSIT6yZgz/gbjJ9Rat2Uza
g1njwEiP2peOPQCk+RRGd7Jq9X0eMJ6GMirsJbxzzTRyfSnNOXswB3uAXxTz8jZh
YgD1c+g/LsDsh3v4LPhB2aDwhG2ldYG5nOa7gd1BqLr+RGDViLFHz4HhNHVK4A07
`protect END_PROTECTED
