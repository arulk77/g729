`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dSi64UNMdZboxQLmTA3JR8YdzT8i8ClkgQhyoLgZIZjvtfS5R9/yA7tw36kStIVA
XM89bkO1taobW1f8J+1Xk8VrMsPR+aYIZ219aRz/iBiIFiBrb4DQE8KGFbsWbowZ
1ZC6ivZUV5BmSHN9P9XQTc+AjkvyUKUNQ2zwNqW72dt1O03e1hwDPDpQU/PvGbp5
V4nSs43PzmMB7cVm08Xp1Lkhuq0F77dXpsWenWwgn8iyz37gvyVt+Y4aL9YRU36q
j52T2r4ZFU4kinYUi5QSVlFg5cnoSII5rPSQn+OgWGbpEkzMpgc0pCPdfbJoG2TW
V9yRm5aECKAnCxRriO5tO+wC398IBtNosY4giuY7Up0=
`protect END_PROTECTED
