`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAfMaEFPt5c2W4OWzT7PcpFqUFvSLHjP82fv3aV64PQgz
W37gnsTWCG8uDlbTiChL/4w9F8ats8cfVWYk5WyBF82gbyFkcx4M4GnEbaYFypHf
mwC+7eZMAcPpIDwj+pyIoCe19kZuKOr6mHFSnxJJDX5/4/8fbO+hrcs8KezH4/UA
O6LzlC4wzIEMObcKU7JUBXbd8YAQzDukmyrXsOAsVixFxQ1Xgl8TrUb/VXcw6l+7
j5KjcXyZBS78DVs/I+1Q28fwP8Ua4pfbkLyYZB4ihj+c7WPp5aK3mBC9rNRGzFqX
AjLRWT/BJy392Jvard/eGrocv+OpGom2MKvUuES/dU/WiikiSOw8Xuq//rwq7ZML
vXKZ6f3kjlcTMkQ9Anjs1cdN4qs7U+1njT4GUJkVQ1F+eMsss3d/9wtuw9z2xMry
y0KZRY8/gVWxNxDc+lkmU0jA3SzSPTuDDPwb8v+Wh81f8w4m4wywCGKGGxmgUC1g
xRd9V7gLR26HiBqLCBK4BrZj8/V3AkZbQH3C2WPrTGcO30rXB/X4c42/3xW1FKq7
RC/EazZH5ohAuEectFo3ocyP1ZKNfkUvJpl4TvwGFqkSFsrxTezw1d9ngG0xV6p4
injjj+j/HNfS/lOOm14e24TVxhxldg8jtk1qI+xzy6f/oJuOqlQhi4/BrYo962mD
14z5Cx+V1SRRxl4ZgZyKcGCjvtkTRMWBfjRI3Rq6Qo/98gO0yY0ufXSy/1a+jMeW
eRR9r8+U+BqGjLo/N7a7AZltSY2wi15g7GVFnw4VuFo=
`protect END_PROTECTED
