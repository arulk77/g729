`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41TKWyo6TiUbfYn2OvdI+7vvuH77gigzvV0agbz1X6Jt
LF6/SJcqP4Y5g3MqfgypHfCfb9QEzWa/KKJxK/bkYG3/bfls4ZCkudhtdG1aAMsq
dMCIxDcqJ+KQ+ADFSAZY5/9B6Rbcb46fuwWFtD3cqj4pcFK1cLCuqA/mMJkrR8dW
uQw7o17v8nRIYa/MlM8wp/W32zk28U+TA81A6b01d/iEglA52OeAI9mpJlchJZu8
YLQ04g7WzB2yca2SnfgFt4t6ruXMiceqOyutFsU1LWvUQW1zi4iiQbVZ9cc0iFyY
3hbj8sXpUVmM/rtRg/YxSw==
`protect END_PROTECTED
