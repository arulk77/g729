`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu407nil9vHZXAvkWqXOY5U1/e9E8a2DUmo71typIHb9TE
Y00vo27ocqRZZEduRaR/sIODEvlxrfJETwX1fQZNY0vWyFvkKrmR4dbgS+pn4wtW
3/I8EIeuAyoiOPF0JJ7ZCYoawS0ermgDa7Hhsc+cUwY4tUuQvSQQrn97Xcwx8sB5
FOrV4jD9fcatThoxtRgKnpRBixtPxZAxQ18Jo9bLpIXESOPXWRk0a2hg0TpMPEe+
w9dLisfxjNEE4n9jcrPV9o1/RRJumnvkAhYo9vFc2EUfWJHL9PLvAj3f4Su3WVvk
iDcX/Ydid5syBr7YJb8mDtGGZA9i77iYmRLcUdJ5WCdzOET7GznnEL1GbQpoZnMU
1NU1ixooDSkxFhtOJBGBVcDtjod0XaU3SH7vfpHiKmyorMfmKcHhvLQNgewEQ1rk
ZyiYZ4hNyjIgUcEv5HQuUQ==
`protect END_PROTECTED
