`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48Zt54cqRVy4k7KZtfYzzFm0YDnKq/Rk85DVIORwt2P5
jSxVn+7dhgTpqrqm37wqbkQF84RJnAydzqIbBJuSK1FsdxUzrIXGxrgTo5RV4XKz
3Bo9hiFFnlRUDc+hdVv20kaZ3h72qptjqAsk2sfubt5aFQR8phIVA2CBx/kt4nY5
38wRoinMhhZwJUwapZbFJEJ01rJ9rIaAC+6K+Bcl2Fw=
`protect END_PROTECTED
