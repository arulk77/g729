`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAIJs7ScqKCQ++RZzQLUrvhAcef7TMUfMbMxS+sOhqpz
D+X6Z7uoINEsgP3vnpkrntB9+y6UPBQBaNcFJpWXrA0aiTmhhjHHPBrzJ+Pa7aaE
kpLA3ZBn40GTng9Tzao+VLyyNasvRa+46v/1OkppCFnGn5Fr86Bd7a2uxJDIKqH6
SzxUwcWvul0ypElxZURGCWSPC900BrO4vxZBFX89ZdAwYD47C3viDFCL8r3tI2Uz
dqarf0XXpqRwYlZKIdqfoOKlkxq/6YEpEQb/E2tB15GCdqpXxnT8PuX8GmclnvD9
2Oghf9LudnA88D+ZMle5yqaC4Vtc2Oz+UxSdy2kWOBYbDqg3UIBsH4TsPa9rnAwM
SF3AUf8AtvRfNaWNwjaSfvOvA0Bakih8tOBVN52G2xCEtY6WTkVU7anjWr94sxae
h3BkQykgPaFwK+CVzQPW2SY7zbQx/dHPIKv41BVd9EmkdtmodmqRmTWNvHKty9YK
3THBQRETIS7OvIhUwjAOGJOV/DRKFCCwssPGNYE8x1Ls0vDSetzQdYP9hYoHO4YU
Aoy8Q4thZdVP2oDdDWJypLNcEREVdfvl0EegQKDL8g3O7tkeMGmJKVOwAPnK7enr
vzaqQnYnoFekkIw4iDb48WB8SPavy780JwOlASbMF98OpLqsRN7kJm6/9UmQJ+At
`protect END_PROTECTED
