`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abEx5IXDnxlC5Q5wNjaFSu/kNQdTF/Kea+VB4+BCZW4d
iuLj8YJ0gRFRHHceegTflkrR7I/prUPjvNHGokBvn0yN1cN7a8QTKmC6SyOTilug
Wu7hoV1s8oRf3xMsT8+eVJluBbK+IFSZjmjdBbS8hpuIlvNiL4aqLT3XhCNthNYu
NWdWbPSQsv3+/b6ObJOkdSUNhOwFf5IAZOTX4aqoS4f+xiSHJDizHKu4rse6JCiQ
3gs3W28as5Ds1s85hZyvWdJPJZrMOC/OU7xGt/RFN12OXBh1+RVBN+lGeAGU48nb
OL/bE9H1YAwwiA2OChiswQLOGg8SJoCdYboEEcDQpoMFcpzE6G2yuKLKPZRHt31u
j8O4KIhRgeaPFu0YpAjhsDQvZ5yes9K14DLGpOm7BVdsspY1/lqeZRqrCoeZl3Aq
agYvl46lunPMSbb/f3LpPANzfOSc025LA1JibraIRPDHRIIYt7ZLneiV9geefQXq
e7z9kSwbDz3lSrO1SsLh66Xl+D/LCytBgI5iz1/eil7+HGhJnpWI4hVBBz2MYQh9
nrCz9u5LsRHOTU8Wa1T09mTK9WC3N6Qf35QHKKSdTmh171miEQKtiU18n4waHqaZ
hcTvI4lebdrMN4ZS7QP+dWsplga2PsVriMOZnIiuY7gIELZyENmrLGd+J7kX4Ajh
vvto9XsvUO+4p5Iv8kiqtG08G+DjsXhFNEknPyLSEHBeKmibOGDS4DYlPdwXYf8i
LF2jDcy2UZS1WTvlcGzPj6id2QH+azboRBC6Yhxo/IhkN+MYHU/UQQ5Bt6yFVDbM
ri/4Bd7ALjKYEJi3fnb2FbJrKqW6dvQIYgAd/ySVfMGIwOEXZVBvHUE3D45QzTef
EpIdhrghAETtDedfNuizsXFmIQf1IqK0vxsQbTAHtwI=
`protect END_PROTECTED
