`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAdE4bErkXROsuBbTnIQJIyR/AbLLOFWUpbwRfr8ZuMob
zNhRAIlMFBQCnSj1nRUKgS0uA92QQc+/RDLyKAl1w5rZO+jM34wKpqOBRm8k9Rzq
FRK9/K4x2DJFuYuSuc+q6CeHS1UnoopvB3mnF7gRu7k/ItGD1TQMsT7mQZeBEUag
bn6oXMcWmLaaIEOPFk9t36MDad8Sfce3HnnburE4FiJDzl2djkBmCF18gbm89VtK
tE8kfsaXerGmgV6ACp+xyue9i+2j6vZcahgOzcIYMMDnFVjx3YcydH75lZOTZn+h
hKIBOVCciOVVU6JMgdX9RyeFjwZ3SuFqa3MctNQnjRgyW1mxgQO/Wc5IUBGlzkUX
S/GeueYKyGeStj0c6jI7jWlM5XLUhQJzuL1MMLdikIMdjXAdLdMei3XlYrfWgB/4
AomBGomhShv01U/mGzizMN3iEuiVyUOyef6gYWQPq1HWQYLdcY8ZK9MqI0soHYj+
vXtFKFYPMG88AujQ6J+5YgliPVfX8RIl1mF9GL6gK0DGB0XLYC54y0QqPCYdihBA
R99eqsro04YzB/0qHN2XVe9sP31Vkb77oUJ713dDVu/slbjDHQgJD/hYJzRsWO26
k+/6xsrowt1oPXGXaQffeZ1KLEoEx1LTSWC0Y5oz44ZjcYotNZsVYveokiOu/Fef
1Ajmp0tJtqavGNSBzaxRKFPenRGQUIHsHFtc7mPZDPpcBFHJNqp82CNVKdBW+WpR
9cFPRKIX+LCUJHI7cl+Ls8U6T4De9QngAyxVzjq9s9KGKkJ/UCHzCuuoiVk/1pqE
cE34oioe65ErPlkgIuNnMxAHOIsXgLPJrlcseQ/HDDTKIYY1KME17nwk1K1qm9tk
fn6JJkkLJB6TLfd7ebMnFw4OjwFAQN615ddIPKWGsM20nq+jHYh6NYIU5Ja+GcjO
mCJSD5ax8VlKGBK9WuoKrgdTqGjOsn4zyp3KuL7v3oUcx04DCnyeqOT5eDpPaSbt
FlZRIcy4s8ZKarynhexnzAmuyVXfc8Tt/JiB3tKdg3dtDyJjSO3bSlnMke7BtAyh
g/CziBPYsBdX+AjlmMFm6xBxe4tRN3LQD/beD4S19X/NjCrQAu5zYt4QbeYSpDHq
xW9qbZmfvkkOzYnwM+tV8EMxkd56PeeS4xVLOBISZvNpXi9pDFcMgFF/9Db7hzpz
KTIJv1dO+WCy2X4kTMzSB8W+AT7zS/UF3zuK3DAj74R0qwKAOAoQ561XfTuSRPCh
IFBK5eY16CSYXfH2Gb43k7a/7pnufmOASqgVYdy8BxNecVGfUq1mUuB+zUf/WHJ7
UulE4n/aUoPnzKDeE4nNe4tLSPdMCz0fB/VqygnyIWAmfgjvX9B+V+BMsbUkWTHR
6v7HV49rod6xiwaaAoDFTHAhS3nx+YzSKyiW2bzqxbgav+PYD3OHbP+bEK0L5ohJ
rWo7ULWsJVEDbhc7v5f0t7sMNXy+GCVWQhgLGmTqNQR5k9zSY68ysJn9rbYvUOiz
GHIzv/KuEmFHsI/iNW5U7azx8emB2aNLyXcQX5AkmGqhwb9weGMjm6B3A2e7QxMK
TYiqS1dTCY5CEkftWQUxkqoq8JXiQiPclAvj/HGHxw957osukiFKIUWVKyKfrq2N
wPHifkRqNpOsqW5OqC61/l37MEiOlAQx/KhcO1U65TeivfFCVmHl1CZysujX4fCL
2ZoZLA3p19x/t1VD5EaSpyBOV6gLwvmn6ePYcQGXrcBvhu698N1ZS3e8ZwEJpz7i
yDERs51dpqEuosaNmN3dm5B0hmMvJ6i3Rg8B3fMWH/KsBccpkMwa8oo/XKjldCSp
`protect END_PROTECTED
