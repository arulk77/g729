`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLGZGFcHjpH7MChCCqO24gbIUonKOB3QrTyNNs6pISWz
Ce4N4m+5RqqxNZBqt47vidY5oqN2h2UOEco6lAeQ8Ja5oiIstN7m2R33p36Tha4A
dFTKxarO+d4a2Dx0yOqi7zei3ySKqz4WtansXMKSXleGuDQy6LeBO0mYnKRWC0AF
8kQlOXQLCzY3JMVk8gZ6wj3vHEYHurhR4T0RlV72mYJczAMafv1VH4jw4UBr8/sl
rQw2R/8d9qdYG2WRTziM4suherknfwzNbHVf9Ob+Tz50GI97YcvJ1P3ssxEXkbBS
dx/hCSU2QMzg1P3RcucPGrrRz+i1rBEGopw3dAnMpf0=
`protect END_PROTECTED
