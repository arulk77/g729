`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44UeTNGNYY2f+5Lc9FOXj2OIr86dAzsi2hXxwBMTKaAA
DE70n/+JbQf4+iP16iEuu4ecPzhP+ngSkjL4S033sg1Jsqa/KEzfGltgO9yHGThc
QigoeF04ed49nAUDODRRwewKH4I1+Cw3LsOryo+sljNpLNBxjMuCFj+mDjwi8lUw
NTt6P1rfdOK3votT2uessQlYVX/hC6+KzZTsdeVmJ0GMizT5vLe9vJl35Us8CGH2
YIuSreUzDQbVoW1Dxgw3wANLu+HjVDp1Endh4OIMyNOl3IhQF9bVfzO3wlo0yTy0
rzr6DvvFunWmFZZM+pZeyg==
`protect END_PROTECTED
