`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xXWe0x82WDX/dKqM/EjC98X0pIAhQO9fL4+g+o+pnkg
MnhXhdfyDWhPdLRo587j7xTxZ/vrHKx+tktWPmFjTOpaPsm+8l/q8Sszt8PPG+Lh
dOefeOc8VnfyKIYtS2OkiVFiuAT87/vMfhTuq3PY1FSePRdNduOl77V+HiNSE3KJ
waiy4Ck471exkGQCFXKliE07AO7LldDGb10axZju4O8XTvHEZehSEsJWhB2uyqrp
u1RjDS2DaF5DY5IYeHhoVaaX8JdZOP+wBaOn6sWi0BL+5tv1JpF1WhkXnDjd2YKK
v2jzZuh+jK5zID/eS/Pr2WRLo8JNpUcG3IQwH+VjWmzCMXOg+I8a72zyrCj1a45f
qla8UmdHHcJYUVUy6QNeww==
`protect END_PROTECTED
