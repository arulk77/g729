`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nne1Xj7qYUoMJ6ULXb1ly8t0O1L5I51a6y+ndGUmYqMSC+2faXHNmwAbk72jT58m
e/bIcjrg2PH7vXG3O9cuji9jfRkcnCLr+z10AiFq+UiYjOCSI4IxYDYymzKt8wyx
32kHPOXQIOIgT7Ci+HfcmsrkGNVeoe7qrvzo2j6K+Z5WiVYrYxid5NjteEI6gzCC
apoxd2UeKGJgQO14qJkijydSFtY5b8gCJv5FXT2e2OSAOdtYwZdxKt8zcJEVPtij
w+HvYP6QJAz5kZyQ/UkZwHslqBWbsOCtxXkpHdCO1odnY5oshgFo/Jq7X7p1q6dz
ZsYCOCvE0I6HEm0lKcoH/fUI7NlmVWE+P+D7ejBS3BG3e42hmb0hngBTC5xn298p
4P+jncu/h8Qgqq06QkW9eruOhuuDNQ44+8ZUx7F6i6/1QBF+AafFpDXaUVchowYq
8Sz82sS/t6WWbWUvKZhScG8E/5LfEpkpIYt6n4yanteRC4D580DEMw7gu1imYnHw
UTk1Txk/TDX4MsdgOdijZDLDpw46AIokV3+OmhVe9IySsdcmY81cttrQrdKrbPsW
s2oPBWi5OrzSmjY6sns2BadkeXKNBKL8oUr448dr5XgwUm4kj323zbvhVvdE+FBk
Gvv7f60Bvv+enJ4foVEu5TRZyKNB2KJcwBuTbJHbmOS4Nau49bVw3p5Qdq5U8FXi
N/kv/RAVon8Abq3drQAaw6X56LNhuMvzbw24IlQEDYgu2BasEWcuSBq0t9Dk5pC3
IzAkIF8afQu+RExutjDtChzglxBdqkSEHCVvgwsZwsXmnTQt51lFfjGjf3Nff9Hp
sSwZ4+eyoSoNLZssKB4UafyV/TEqzBKdTSzH0uv3y4RXbN2WgmVMhcGvRJ1pVasy
C4ZzAed+xJLDNQU0FBHjo59MijgPwkdDbRPWxglEwW5EVsVOnx9p7hZUGS18wJTO
oxXRgv4DiJIzlQDMTAZueJKptSMTI9I+e3OR6k2XMqzwXBxp3BLvqLcpK3Pq3irh
1yPc2dQzKl4lbJ+VKYZRtBi1sULldSypU8V153xkFspBrd/vjZkK4GCPc6JR4Zkg
r0MtCmUtRfdFBQ50gbJx3WkyJItJ9VaKY1CanHHHfw4DfePwZ0NxyeJybBmq46m5
fRywZcBcnSGioCSw99jhHYmbdsd1bzOuOfNAZxd5z45XQLFVXA1/5LX6bstrUfx4
zKp0QXty7P9YuTmhqv3qCX6G77vpChOznGcH0TaviQITOIijm7kTT+sOnvlKeuDD
FssteksYNCGjEEmDh234SJsL9eSZBDKweCNPW2XKWNovNJXYG5TAh75ZiEh1H2Zz
DjjHakY7tSlaAzDsD6gCtqWFGYJLOGiCL3gE+GWGqEo=
`protect END_PROTECTED
