`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC0HwTtlb862pofreUJCpTgsxsE/1vsHxzv2XiBT+8ut
53IovPDyZiLBZai0a9xjaZ5CKxFwcnppHMmTubNxGKB2Es1qBDUNLBvrWVTPjgRv
lCAf/9I4XchaoFuj2aOD2ukv9XwqJkf089uq1C7vOaWAoVwz0LS/ELogQsZjJVUx
Th5zSm72rLN9PrD5976Yj5DshiF0qB8qqOXx4E1aldkaF9z7+KgSVs6XqH+1Pz+3
4NYENapOf2itHnQCFLpRUR2jiDt4pfmAetCZGZn+W+47K5+7E/uVCAJyKH5ZFR1/
6JpCJA6orwCwMAxwiCOV7YMPtZSzPS6qM+vFcZJxsEPRV0hBErZN+9OiBxRHEHZc
`protect END_PROTECTED
