`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGRE6t88Sk0lM1GsZNV/V5yFJGRMBNNzZDlAVoLA12dv
SXhUehWVsNEk2kEbC8/aZJuQj7NfuC6GK2OZlU1JlzxLX8BkXys+UnAaHMtr//mi
h9qCTLZLJ6FDJT0q6rRz+E7bSJ6jlw5zPWcOK/jrxASiAyUUuKf4sLqVEfoU6D0c
JcJ5i7TaLlkuo4+wCBKuJg==
`protect END_PROTECTED
