`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu452DUnTljsZpc5iZ1EgJmPor5qFFyklAcFqFRr+ZYh+u
JCHUyEtJjdZ2Np3B5YI/QnsbAj4EE444uRxr4+3AFFeRMc1QCCUat5nvdR3dyKj4
iWQBPdBRcTnixudkr25i+ql5du8PPxm1JTAsHxIRwFQ16KJ3C21NgQ+o0uv1Uh3N
xT7SkiHxs5Cf/HYJkrlohsWsLb3tK7m0I7aa/j7E7UQMqLlGwzM6CtNMQtpc9oV9
cVfBu4tL09KIDUAOfrTfYu8K/G7duUZot2PjZ+kOBjyMW81jayhhWhsv1os2RxZi
zXblBwgIDvt9Hx5dYFXzDA==
`protect END_PROTECTED
