`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42bF3Yld7QdKJe2IEe2B0QQm0mWx6r464E2EWCspmo4b
MPxZdn9Cq30OI7I0NkFMJItGOTDUIunJSVUXl3DGBwT+dcOPlvRpBj5uGZTvgDIv
Ev72PjkTSu7EZl5dwt9RKWTUTUHHZOGn87MkHE5oTF+TQA3LQZltrS0UaJA3cO5e
EtnUIqwMkmABMjhrP1gTvEOXa/LASCS5zZXTjAeP37QbWtcqB26QL3WYEns8sj6v
+v8r/IOpo+XVNuFjm0O0xFOWk5Dd4VCFzNTcRQIf4Xaut/SqxsgUMVdcz+o3rX0P
71HO1iSuSgHWFQCknYxDvo6UTrgfdjRKtJxBPjBBtaN5wrMy2zhHtsJItv/xdAa0
HLWf0Qsc5FTlNbnck+ccRCH/x//xLRltZtAzBAx3zfuJm1y5sxPuTzrhffDIGRU0
pIXJ6ApKzva3QxCXSfb4EsNA/+w+8G6jBK0o3zi1Hz1KTXEpgvBEF6Q4Z6eVGwEE
`protect END_PROTECTED
