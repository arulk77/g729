`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLcAKRr1IxSOg9aNY3+Pvr2wFxJ8QLgnb49YlSdGLmc5
Mm+BGYn+p3IRfNPI4lJ3xvEhKJLy9j8pJNXC5wSuNl1hjvAV9RVrTSVjYmhJSt0g
GEW660gQhG+Yb9VtqFP2Zghs8tHoyfyX+TRDXBnGTi+tYubNpDWmQlq6C10pD1H3
CuX8ZwSyIcEdlCUyCpvWonEAN6r+Ch842RnL4nG4ueJDFOZG8U8MynOdEUZshkcK
`protect END_PROTECTED
