`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xoArcJ8m9nh9Eb9zR5JPyfTqmCdeju2EhiAHkC4wtj8G1Y9JIy1ebrIXZVO9aQ4J
WDhjJxJBy/wmWlfrmK3EeCRZ+LtAUalHv667V460WAcq6vdU6S0ZbLC/ySUzcmp3
aP7e2LR4ZoR49Y4QgkYKVU/nNu8zxFOIG4dfgAhvXDcSiEfV+GOSknrb4IQfcTyH
O/FAmzwzdSzawhAazLsVLjeII6PiHsb2/iD/hG67pi5WLNiNITCE9O4y4m87tm1w
+Bx/zj+Dp1iw94LMDelAWinBDYv1iQOCGizM1+TgLw8GvkG/6z3Pcg+ECI2N2oU6
YRPSE1wRyja1iRhcATjt9i97ChOUh33JG9t29zuTY8I=
`protect END_PROTECTED
