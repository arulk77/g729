`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAVPPJY4h6k7gI8JHm5RjGxkJpK84/qrk8cPTgV3/ZSuv
GBRFdeWaR0c225QEs0wqZ0NdQOUsYdjcfxLdGkOyHdq6uaccb89kRQrTxBDZw00M
OQpoIDu5LBstcgVlUVFdrIGh8Of7g+TnBgG1BfFUoUNy1WVUbstrSBxwM11OhaUs
XZrA5GfJfxZvRo3MAOS34pam6tyigWQ65PeNWNhSN+kkelzWkkV1NtEv4cBt/FeS
UQjoCMHx+NW2nWjEyoieZdrd5GIZKig9jWMPi8TX+lyVAH24PA0b9/Rcd54JMiFb
IZdPKGbbptrn2I9pKP3fllEMA7fvbRQT0kZHbbIaLIusOJm4jeP4gXJ2zGxyps29
5C3kFEoNJIwZeNnQ+V2ZYIJwqa9WdIGcUPZrFcOY+8t7Rr5ZYkeUR6GjNHfDeUvc
TbeOW3D3Vgda3Bhgk3L0LHxtsTMfAJJwTXO4xGhKJHHAYXJiecaK/GjEt7Bm5QUw
goqvjP6aILLWFusvTje52OOu3q011CFZCUw+Cf1yokw6R3viKlzy0Yhwea6yFzio
Im0llmXTtKR0LXdrQvB4SD+7MRI6RBtyAZh29ELDno1ny54a94uX836CQPAoPDEW
lJ1U06ga+S1gDR4WOvhSz1EAfLgKcdhiAgzd3w0/92mX+Gh0l8Q+nBSoJG/W0wOj
tNdEfzAGxQh5XpBU9ovgx0M5jaf7aKt7R9e22To6mF5aDCM0Cyan5mlkQzJ58nu0
0dLeDsbbzOPIldeNOTnIsw==
`protect END_PROTECTED
