`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHNFlVA/GG5Jx2RlGjvE68rlIq7PymJEX6Jh/9sNEesX
/1QqvKcEJ53tUPutQ16GwWoXO7tB9uF7v5BEvgmGu4x3Mtl+O/PWXuVFVgg0PI+O
CHM79SJCXZZuBesThegZPXwEMlyQ5Nh2RwZIqiyjpuOCA/rYdffV4SLythJY09XL
z6dhe8XlAjrau+5mlhTOLUBvz0lcgUJQrz9nrS3zR9LP1EPMGyoYr10+Stxq9v+S
gJskSErWtIQ5N17GeS8CyN4qdAYidkg08EyT2AEV3YPmIkaWaBHe8/tt0EzEY5M8
1WUPuaE/bli+YYFr8ionHw==
`protect END_PROTECTED
