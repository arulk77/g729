`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZXWdUm57JTZEnjktDJAOvA86CPeBf+LH1hXAwrz9Gn6eesiKl4vSDu5xY73NARmG
mCFhuqf3nJsS3urd7d3EQYV4mlT8KjhRI7gc8a/O0uTUcPBe03UwjbrXHmFhSR0f
Qyk3RsaL7bffOXk2tRYRTFHnJuXbcPKeAGl0E1RPobhNdptv4laHzTf/7Ia0gpO4
+03fRzMUa85YeB0iEZSRIM92nUCLtxsRLcEiZHn/rWCsbEcZv8Z4Ij2cjE2yMxwe
3NOIdtyp2h7rSb1vnbgMS3Cc96+WIfDjiUR4pepCExA=
`protect END_PROTECTED
