`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cOLkOnM/bitqt2OVdapdTT0DGIzHtqPdPaP4/vCQRcGi
DDTF84KyM5hQwKGK15bD6Gz76vmwoYgz/VNr00NrcQQyDu408mB5Veg4Y/Yv9ptd
94jEnhR3N6KloDB/Es7Qx/ZzvMUkgIW9TWMfTzCraeJ+TCAa3452cwWUqqmzjHaL
`protect END_PROTECTED
