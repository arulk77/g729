`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH1VEh7EaYC1hINod/wamaorVS8zxr/w7AMnga7Z3125
2fXUQpUh4cUfC4kPzxwPQ6kp3vEwQ6yA7He4qZ5wW9OmCOQZuphqanjliJJdLGlg
yoHnFqhuNlaNiRBQrZ/JN3o6nhGLuVJUr9GQK4ORjnlmHmSvMdjV59b8U8o0RSHo
IldaP0WqwKOpxKidxBHkPw==
`protect END_PROTECTED
