`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveALyzXmLSd8SlpGFaAZEGFBSo79ibDrAmuYnovnDLmZm
T63HExgfTzGj0JzdNseLZ+SAPxfsajqoyyL8F7hG/Lk3Tg/hL78b1hk3uM6kclGE
716t+/mzJJyiZRSzWqcP8ztvcRwOWSFVLetNv9KT06/3kJ6TaIWUoLiB1bGchoz9
`protect END_PROTECTED
