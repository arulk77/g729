`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAheb9cnbbi3PFvYl2YKTO8k7QHeESGHlyRfIVzpCKP6
tTOATpYRRc9fTaCg2kywSffG6lH+hTNGWr6C7FawjAArapr/ZlsMBZ72E7ESHBeY
YYmpRGtjz8eCVJa1eo6kdxRQZjBDkANYd5kE/IvXsIH6dG4AZs2oXuhwVii6m6Q4
Z7yJGKOxMVGouXPrIeqOYgfNCcaHxNZ9olGzuwuMdzNmUDI+00Ikuvz3VWB/PuoX
nTHeDTOYryB3fpl0cbpETclvsB2bRq2FVAPnGHGS92fyUBZeeHa7f6WmcLRvN9A0
E9rWQvf8urd4m279wlNIsbt6E2KZh3PKyTc3SguVmA0/nQGGTNR6oDVBPsGfwTse
YgPhBbS6tHUGtxVt8R/2Jw==
`protect END_PROTECTED
