`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAVFX+HKc4s2Whw2/HqE11Re/h4NaN2Dl1kZeCLy/dPG5
nP+pUqwLiU0SY/db9IjbXr4XvrvIqNarAUp8woip1gFS+JJg0scXynkpzAce1Nys
fPii5w0Ts4D0iMoBWt8KAli5PRIfrmr4Gt4dHBUFQNNZhlLSAKzHJN+kQWmr6aVg
nzqSuMS+KoUxDvLxgIkpA5N/VE7FCR8bQxhsCvrlgHpOKrMab6caCN4nMF9cyZqc
ROm9iZR9Yj2+lttzX6jznkXq5BvqraQWvPwkUmlyOGJdBY7IjfZCZzdGbkVifqBV
DBo1D0/iNktr1gn2bCqjN7TL1J3rDWFX8hiWVJuayq1pDB4N2akz41tZLA8xLJdx
szI6q1c/+cBPj59FC15aVrGHIhWrsVN5yTiHfb0qcXX5FDH0qSLKMaCw3OiHON+m
VJpckPB4al2g90zEADxh1LNRzJ8Sgu5ySYHRT+U/OdUZACcr9CMEisAxSBCdmSEl
yFyqMggLLDpl8XJ/duchJqxn0fvDbFsCA6ujtifpbn453rhLSResqLvvptEw1Da7
mYSAdFnYoSPvDjrdDN8wySJl6e2EQn7odiV11+z+1k5HNduhYLfTJnCiaaXaMW3q
8skhtAF1lEu6HPoEFFg+ZCNZM3b7qxwOL0eukHKqEEa/R/V4ugRZq95mitUQp1c3
F98zMX2IiTW9BFpR+7d6o9iNk9dw1d2mvTQKJymiP/QRz+V8p12uHaST6OfAm4rg
FItW9YP1Ptodbhwnbs/WdqkQClWxW2I0iGQn0Gk6R9K8j2DqVc2dp3sauhwmVBzB
L3fqYHLJMM63znqfi5hpvWOBI7jSCbYiPJlv7xPpET1a2bjD16nKnZOgovD+gRDU
JbZ46bndCW86vzXDAso+OjXRQl/m9vTqo9vFBpr9ozSG7d9l8N1FgRBJ3S23uVwx
MjhSqPYjX7BS4JVOEh5+K8FoAbS+sfXodVujjJo/Hh6mbIw41G5AHv6WQBE/MMBI
wE7Q/vpWdFykTmGekIzpdDMzV0RIysSurKE8ZUD3VuxRKGDaPWkSczaqxtKRAh3Y
kxgR5NK/caUBBZ/n2Xm8hl6yssgmPHUGmmHTJAyKoV8Xo407PlAacO0MrXWCkL29
LfSDuHQr5th1ZI+Dr7Px6S6bVL5g2IZ3cGT/nrPGb/DXxAx7nFER5x+Qn2i5WNc0
VyRK6NeBoh5HBZZPiKklVaStSaFd0DZdbRWOzpNa/b/11I9bY8XOZkq5jhJmllwJ
lLtLxfW1MGyxsrXQjRdgdPR74Gpt4DrETzWRolJVKdXqlB4Vh65ZHbNCTmIxBwyq
ykqf+FTmUpfBzGotKvH7vOzRHX+JzceUTa/YGgyg+iiaFCx4M22rPkzJyud87WBU
fHSyamAV35Xzffrx7Asjs5gaX4METSqM1HaTjAq41Jj+OZAPhLlMo51kMLWLZuqa
f+C7TwFMFNWZNc67gy6QeHGouMvL/gqMDm+t6DaNKLEGaz0EVnlcBabzdwiFCNWP
4FDJWP2Xp1zSthOg3hnDnunW/YpfG7EvarlgoNJIUQU=
`protect END_PROTECTED
