`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN1kqkY1rrj8nlfgoyNvQERRb5lJqcFS/7L1hVb+ToRFv
J7liWsZrPZD1xPt6NyQG1MAsDwf3p6LQAAjSZ79sabrFWIih+x3Nkp2FC2CfTt4r
NAfs9P3NrE3If3iksAMeZsOxO6nG4gwNVkrMTyRT0siA9QVrXL2DhvkyFIdQ0kOB
ftuienH1r73q48JbenJkzrhzvQow+/NkrjL1AdpQeRxx092/WM/LfmihrZ3AxgSB
lLg4q9clPwOZmKYk7vLrJigjhag1qCRNjiCnZ/hx+bEEDWwyPhA8DmenhtzmaQrk
lm2Ozcd1TmbS4/xwgONML1dfc7hKRwmNx4E1NNrH7uKeolQM4haiQl1BEEh+I7i3
prkzXMIfD528WMIcTNW47yKOy6RdhnsPn2rd4u9VmGRSrNmG9qxKrlTA9NTYuG56
FhdbHav3aga1KGuMKDLBHz4BUGlbXfaYcPPswW8njzV67kpIOiowI+NLVeKQmdBU
QIIX8HitTMMqRRNr5vKb9o/ZbKmZBvy9WwlfXmqk8+DXv8qLd2rloJ7DYao4AjBx
PXH8wgK2CfwxvCs/HI26Kqc11Yv/lmf9vtZzxIoQ8RFNiZmC53CFUN7cLp5B+L3S
o2TjQFdHcv7v7Lr0Q3i6PL3UNAJdMnr05qV4yKHPRBKgbi4dgsTPzXvn3BlhGusj
Ro/Rqn5A5oWz4hHOJcj1pKmItbjaBa52Y9Od6NbCiu3JpqbOS4Kg3Yc+WE2sslNw
K5Zb/15Bl351vx7Jywb+HJ66VuBVMWZzPPzhHXQFzEIL6KL/l7F2hBhXH17hOHXa
nJirkgexiM0MKXBTeHtpkRsqftGugntiL4AmGfXEnws+u8nKVX/+8ZfZnp7veXIM
oCOaHE0T//csIHT9JxzhZarckLt2Y9rR75mJSbGaaTQAE9Pn3SO3CJJacrU+ALS0
+2rB5ywYgv4lNqxX5GqXbM81aRobbj6y2Z4GfmU0qAIjMzj+wmlYTSEKHPx0mWHr
m33MKATRxmk/DSNQ2eogByro5K8OTZ8+vrWPbeiGiirJannpkB7/caqyk+GPHrKy
zKvIWJZaf8X411YNC/MdutpfwKapDna9B+FzKyUnXcjMLTUiohDA2MZoGS1GgR3n
dBLNOKYHzEl5GdPPpi05shdDz6e7xFruZk6NfooB2vo64u274ITv5ZoH7CiyPf8n
aR1/XHCP6ubFX3N/TpQ37uB3JRNVSDDF+NckMp2Wfcsq/s71hs/mBf81V2xgS4aR
bHbgSjDWgSo47Jk2tyAoY29+PfsW1+wyOodS6D7DRijsWx7KTUsjL40V1UvmKh4Q
3GVo4hVFjRotTjv5f1bTYfUe5srQBZ5z9+1tNdDxV3z1PZCqlPpUUDFxLMFKxN9A
9aBLUi9eXRERFfJUQkEwvnz5ULPrzLPXgMqTaQH1dgsKQ0TSb4rnvXyuU6NpsY9C
MlUsY3FvMQHcBWQfvsT1aUSbpVDZdUkMwDQS/aVFSI0lTSTjHqJw05REtO8Y5pr7
49R0GVwlD6oH+XtGVrcr1/FHKVWx0ArOu1b4xfadimcnqU+nnjiI0w6hdFe9gReg
oV9pVeR37ui4juxQQCAOu3B8S39sANVU3apNcnjhKeoVwKzBBBEPA1y4GTQJgKt+
1Dx5adEpkt1Itnar7K8W5G2ycM9TfM0svELpSwjaK004pvK8mI4/uEb7sKga1lQb
yAWpaMkeXmKEtcTx25JqITfaARE+Qvd4ISOuVvIeRHlagnYhKH6zgLLaoyFWSYpt
rEvjpk+7taOAxD4t9PxLKvKcQjMO/7EHUoz1qX/se6CjEbG3EcK3V68Al/EBwuEl
Wr5zzPTielj5DtzyBRgvqFhtCbSd74E4M9jmu/TwdteumtXNCwRZYuQ67Yax9039
sivIXoveqTXBG4O9MiM4E6HVNKM8pd1oX4+VuNvU3Sk=
`protect END_PROTECTED
