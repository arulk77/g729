`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGJixySlQ/ATk0TXdtx4kSHbzbPjbGOkjoFC9aFUsffI
ebtrtHZIk+1BWsYQZYaHvSDY1qTHW+qrn0OBLC48OQHPY9jCH9jjy0lGzQfBDu5w
qUogbrBbcKRev2H0QiPcK785XGaLTLnOR9CCb14AZe6VT4bXFFPR2WYs9Gh5gu9p
kNS+WgoZBsPy4JCgB8ANIukB1kHvwmuLngfz8Fn3/kguwitn6Dy68pXlTX3H21VY
rHobXFfzQG3GOtrN/1WaOn/e0zq1e4eVzunXvugUOLom862qeZb309PKHKDjgfDx
JKyJiaahuVEX6W7fgmfBC96J5Y/Q9cTl2lXMIUu0EfCdsb4IIeYQUHJ4ypInQlvw
XnNYJbgdHSOM1rxiE5JSvA==
`protect END_PROTECTED
