`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAeS94gz71uja1SNHaeztq/CiXjvIgT2JGoGfqoiKnqu7
ZW8mb4zcKhn99+tLkZpDTeTXWxmV8UBy4WM3ewfYG141jT3JeOssVjVqwI+AXZH3
UASy/fmMuqbbMpnaqfjZum9ldifhp9rK2RVxwmL80TOMcTrlNzpkBGDvfl49D/eV
jdTEFFEuZVzDOKTRlzBT/vBOC08SftrRkBBXk2l8NwLCkGJEPvwqskkLfj9Gp33k
y2ftDD65pbi8bhQ9yNqQNbx9qIXJqFfRqbbtz6pNyk6u084yqWCodI3A5LPxA+0U
ssRECMftWMMFtv/l+b+e6rcRVemH+IXSwplRrI0xRgRYX9vsW/DxP4GJyICz+uAq
hT0NJ3SVqb1/p8pXMS1ojXbjJBzwaPwo7IY3GAVddzCnhKfCvFu04Gl4vAy2Czee
RYIm6fMks/r70MgWJvjOmvdqRvR5+IkWFWJ1CVl+CxSkRJjhwlGe0pqgnWfv7KDs
8RGrrPsib19XwjtbrJaoRnLobQCc/VrZ9RGrqxh09YNIDKDkoXHs/x9sS5oQA9u7
xvuCy/3cnCIpuBIyJB44aAH9h5bI36vs9rFC9ekz7xjJ8WmTfIFF5M+euQTOTEVN
3gjg8gHETPTGfWgCAEX2UHGs189YYLP6ZIRlvL3YsMhsivL5V4jJh6Cd4rxMEkXE
2dXZoJ6Lq30LZVXdKZ0wF02UJiM31M+AsfX77cXzi/hNPaIlumI4pLawHdU/lODH
F6ljFUxUXhjrNjGCmbmplAzJPtpUBZXEtppMzzBL3NAefMJ0mXgn2Ryzt2Fv5nCa
raziHPlvQObrGlGvPsAO78ia4ocoN7ec3PyQ0jiDsfzZSWZNdAbwcMmzsyzr5VPe
gDw62mXWfxhX3cATkQCI75y4LFv55M21Xo+PdwFHuhj0Qr53LLfyatbjz8rUosGe
izHEMp3px4LWNPF3wgk4a6h8JbXBctej/sQRIi8Qh3a2DDizMtr8pVRUHu/ZWD1H
MImPdmLFuzc1gcFYmIpFlPMey/wqmoiCAmi1TkqRiD64ShNZkIdImLjaFtKn1aNF
DTYlcRQ7YTky5Y8aNppVi0fy3tGlnb9UOzUb6Zs/ZcdeHhQAqFtYaQfi1bDEekTv
ugzlH+cYPV4OoCtOSR9N//QPJloJTy7sq9yFctJGL6VY1+F/8SaDgqB1F75H4iyp
h3mYNF7zwMr/kRBQfGaQZ2lNo1Kk9GwnPRwPETcXW7E/ajDM+AFLGXzv2mWv3W38
DaDrasrsEUcL3mH52iHOvV0c6Ns93mDEMf7hLpVWIVRWwgDMLGJVb+RHMU/5uJxW
XenKvRcJPQQ41V/FTsXSqgRoLnUhi5aRuJs12/yNMEOTwgUnKWZcDIO+18lQ8GC4
4Vts7E79wfBk2FvgMiXITUY0SYbqH0kcW4zT/FCBjB3i8J7Zh/f4sZnTrsKHvbGT
6l6wTpjddLFBvPs3Ok2VkVbNVIRK5dUDfTq7fs1doFQ+69c7hNXiuhKnjILJzXqF
SIjyAG0/jG/CYnbkn3uPrhLvyLSHyvky1qBSwRZsS3ZvY7PxegZ8HHH2A1fZ/iPZ
EWK5fGGmV3rvdWiU49lTikVaaQd2sbQHZgk7Shcn7upsv9EYf87zbPvMweRhwBvf
LbY19lz0LW4/2dks+3LP2w+6NrVWrdIOPPz4bEdutGB0jDxuGdV5IParAboLyO6l
esssX765Z9BGGf4QhdCe+6e+apcbyVH2Fkzgsgh48B+I+2Bb3HWuInh8GYOjdFmP
ZEsTBgoNZXlKKUoQlMBbM2z6VnFiTRLVqhARDwMP6Ectbb8cOiRDIclgd6UominH
geftkva09WgjItACZFz2VCsVPifY/PbrseTpvNfQzdDd88IOzuy+zbC9+IklIsZL
h7kq9O7MzKH56L2SlgR3itkfs/O7/jwdPYmHuY37rbfdoGTmYCV99K2c3i6NVvSP
B2+RTt8erhMmFIloFw7Hu+pQsl0BhE1vdleUluvqF6N90tlbX4l8y5QzGC20puRO
mKVFLjvjTziH9Hn9J01deS4x+8AWX2SM18qYAcx0gPIVwGv72kQTRkCiWxa+B1i8
GdNy1QOVtD7TpBCrODm0UtAo59dEQ9GHsXMc1vynj9AzsdyYduaedUanof5QQ6af
NUmtzFfo8B7zHkZGTx/FNg52W5QLLV39yHWeyP9fYYt8rhvJSkKtH6kxJzefTlaQ
4TsnaPnIMGRUM4iCNhXNJ0ZJ4y7lTlU+ums+UQQIQ7rDILBLN3HphlZwLE8ozoP4
n8uJ2v4Q0b08OIrAv9llZ0kgwG4f4Z/LHM/B9BjJ89knGDrEL8wuZowxxc0Fz1uf
y2KcFfdqktt5HTA9okg+rqrF42pcMUzJPe0cOzrUweiqkgROANnN3q1W36qZ7rdD
FSeinJAaX2wICMxBt1U0YBAo4f3WCpappVCtfqHUYGSqR3fUxUb3YkJrMhlKltFs
taPt1/5YF4gBTTqEmuHeixj6bmD9iOjAcOO63AJ3Epzr0OPvI5Gfk30cL/G78mnl
9uc8w3Pu6hQqRGTR8dytgwdLurM5rsTxW1fq8jSxldAPiNY6l+32F8igkd3Ya7oU
bRpxInj+fOx9AlZ/tliGIZTyvRrJ3D2Y57HaA6Y7QEagZawXyvHCdYzeX9G0/3iM
2+7303pg7sHumQcJiHOrXOtj2CYnpWSrG8bh1hIFCsBsL+y4Rc6nf1aMCunkfX4q
GJpfA2iAqZv72qPKDX5QvhCnav4KbD3lLiis1bIgwm5uZDuhwVwN4qH5p+7+DUvi
dyHyT7iVktSSlu2qFEf+aOtxVIAjxYIKkvRXM92cRXCKmNGdy0/vYLNrJAx3X1Lg
npGe0y4EKfgi/Z8hVMIxlPWUvPZ5Y0q2cVHj6YKxR+bHMj1/GMR+jKlZ5nKZtZQ2
JVG/SRc/JXIz54Kxu6ftIsTu9/cDwhGn6NvVF/LAmMvggXbzMZSw/+/yVfEXtkry
EbWtc/2HbjQYlvd6fIvUKC8sYjCuRiM/q8nqi9j/zVulbYvdvSC4htPYTUSr1O54
A26D/bNo2AwiSGqNDOm6BPD8tXaXvdMHPlRCTAN4EJa+MBrBIHKOpdsTZO6CgHrE
s14zX54beVWzfyqu7ck9puq8oC0dm9lG8V/GYCc6iRY=
`protect END_PROTECTED
