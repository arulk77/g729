`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46GO7l8h6FE6q+z6956amvYH2jlSnd54xgiorKpibAs3
wHD0BDi90wtS3EHx+INHg828buKmZ1AEejcv/sPSx+nQ34SicN4jX+yhfG3uT2CC
aDAQ08QzOTNNJvhV5YRw8JfQBP1jlrOAKy8lPedDA9HKfEBhVFtY72mga5hzHS7Y
jOT7x+XeThdF6ciqa3oUWlNRcZVFmDvc5OEaEHngH68=
`protect END_PROTECTED
