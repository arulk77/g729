`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAQMGZB2dNcNDdu5LKNBUPxa8wZ49Ksgv/MJessAi2uvk
9M4WLASDD4LcJ071ev828Xfy0iHGKDw9CZnlqqktOInoKR7Oeli1L9oaYDiouYvL
1lXafStaDWwyGFIYMUJdP5PfwsYNmqhUP4xddfyCMXrls0bgrdZEMRRCns2LXIri
SgP+wDrYi6HY0Y3ccAVZ5DixscTcvzkwMrXNyPgd2LjdnQrG92qW5xHBbd+UDhZ0
0r7AOcbYB6iYMqTL52l3p9gl1SMLmoUPHEzfMYz+DfZAn61+zXhz3VAlyTUoJxY6
uDWEtvUtuzidn9LRGm/09QT6EjwP0pn5ehnkav1496g5XjwMAeDmqme+oVEKY/FH
wYdAC1kLscr7WA/DwJP7BaZZ6PKy7pp6dWByNYRm5SO7hxD/FxBtbPh9pFtqt8s0
j7RVgnb0utR+LREvBZ1iUdxRXpXNvGXIAHIjixMk2e8eB8/YW+DrwH2CRSK+fjnL
XFjL5BzFJlxXRTboxBadthflYd8QmveE7ubqq5lDZxCHpniVPv0kAATzIxMr+iLI
8S5MUgN5APFKk74sCZKY0/0ICbX/0/8ziI2Yk3zYfPD30ccCFsX3Cll3TpA1KucY
1PKLv7AcR7upP3n+SW3rIVl/03ZUIURdBKbRYB7LDYjmDWa4GL8GiGnt76cgZvfB
UlK3aVHxkRTUjg0QvIPOtFzTiY1h6KcXZz5loci0IxMc2PEFSElx6ugshsCZqFOY
6utvquOe/sag6ZtM/kVgDYx3kVI8A/UmmRaVfYmGEUXjraPBXetBf8Cu4r+SPyRI
bZ2j7kx/ddCy6NbgDvOnYac05A3f98YiCxkwkh6e5Wjo++buHy4IwiYhPE9i9BYr
FYE7rI3lD3lzyMh5mMOL43YZ/0C5U5/MqgrwFXL0XEhRI9htR6ZoeFsqnkzelUoc
VsYG3dKg+gYOtwOt6auD1prV0F6zruAAsIMklzBWgwokHrOfiAI3A9JtTUjbVxJE
6y21XtIqEcP+ZCcum8bPNEwmY8Vw/3ShTQFnsTXQKPY0WTVo84c2qreoft85Lwr9
4duTltrSJ264DpVfOxkUb6S5EDkACVfKPIjc/6/m2oIBXrgDj3IDB6q1MmAukPsP
/Ekuts3WCYQ4aSW/x3Ae6OgieaHmG6n9LLFEu/qCMES40Rr5SykVK+L3gA+bzlSI
fG1txEpF8bN+asF05kaG/ET/BxmYz9pe8AzjfhKVPjXe8/dKeTCr5i9S/bEAq4I5
Bw3Cptad+V16Fi56MLYf1y4A4fJED0CHclWCvu9Y8IEOE/oGg9MObeJzbpAv77VS
JsCTmDTbyQB+BbZHIMTbc5oc199vyxPOpgyDAnTX4enNm9BXH276FQ6d50RVJTdN
FilDTYQ3fqAxWpKiSWeCGQLPi2ssyfQ/SSTkevXiyRhr5RDKeBUGjFZY1odjt6HF
Is14Y9b/dD9inT5VTby7Vq7cbdEE1gSUnlEypZlMDKbkAIeONqFuhBvM+gnn2n1c
cPqvCiRwg30pq9HU7ZJR82GsFqjMHVCeDbi4gYPH9nyMDLN3U0MD5BbaPhUb52Ue
Pzpq9b0MMZyvCTE1t4xHFdkBfh7GkksPG+t2ZNVzCIoplZXmOj8oxhoV9+Iv03b+
bGChIrojKjNdmlv62wGWDMamfkNzm9mYGG9UY9bQUcSOJEl1dcxc/ja2sGg0DnfL
Fmj+5KizevYcXldYk1O4QnwvtAsOmb3JfW8yEAPw4RCaEJN7WOo1/sEFx2h2b9Si
WK5c2fweda2slr2a/fRrmztunFOZJ3+iTAwd+xhTrAjMQHDIUwK5p8RSpMaxr2SG
r6JKPUca8XwKnz9DuLzKbEmm0b/rLksi7sVnkRNpVCaFlNbC1RWHg1qAt97W202A
AcZyj6rpk65YA4u1L1jrdR84KSUQK02ZOnv3DEy+DflBIa8LLBbZf0n+dmOZzZpd
Q6SlrUoqYTlQ/PEfpaIDwZNMdcm4a3ZzDDZEyiqZvpq56xFIqDjadRGURQPD++Ma
sdtKORZcwxZi0pq2hXFev+MouT2SsrMqU7OGZBy2rYEJtq64lY4h6xhUaBwYVwbb
xTCRKyGuPrux4RU4zcfiAYyQ/DiHrsdcro6SdpBHX7nwg8aMDw2Aohfjjt0BlLEh
`protect END_PROTECTED
