`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK48MGwre3mtu6U8ao8AWrf2kwiDmsczk872KNxTkNk/
ZB++GBu2BG5xlOpz9DAWKx5TEeNE7ZnyCbWM3brPPnmwBL6Zk66LoiaL5uH7Cu8p
VNhQd9aM4siYeIvfAqrnr7ht/T5DG9idMB0PCSY/BLc4qejmTExlXKHaKz/AugLv
eMYjKokgNjMSUPGszFRaTbj2MZuofOS8BMrJKsV3MEZ21qhrWv8OqnxdB1i+3czM
W+QIGy9qd0DBJ/Axvizu8TJRWCAFX1gHKi/N32wVrwenD+Gl6c07yZJWNVXGN+/R
ycZKYAD+HvIPu1SXEUOgT0swj8fHFlsJEm/OIGbdW2JhHuUHI/yNrxg3VBPlGr7L
J+tp8hwgB44H462kmURh8lUj2kAK5AtPheFfhI0+NZehkMIpOoAl1m+K+U/qk2xD
`protect END_PROTECTED
