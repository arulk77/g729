`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9avVOGSKeHN2UCtOM4p8pA3E1J/aENQPYJxZNczs1b8kUg0SlFvpRiUT3E53FOhq
O/aLV3Xrf+0AzVGdUvcePce5Ref3b0wiJPy/91K7skKoeY9+mtgFWAdt5tZtI1x4
TcNwP9gO4Q7rnF/whiBBQWQMBQIgivFVR5ioIU5J6ZdWrqy8PXMW/ZixM57ug/Ba
1gjh2Bn6Yj8Jk5JKfVADnXVHPcQlADIeZhhT/FJW5KsaZB7n2aQ6BLBgpRhjBEJi
QwCxJr014By7sqkc28RYd8B2pMuGDThM+43bJrlYz7x6cjmcLL+KJPmeY/wCsGbj
FpkbeMxZpD9A9RiXRSMEAjUbu6aN840xFuUBLm3WVGKmwygxDzTHeticz5Cy0BYj
qzI0aQb4fpntieaViXRxRyjrxNnqabi494Tu5/lzMr4=
`protect END_PROTECTED
