`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEPXo0i8g9uJ+9eu/J9h1486veqAqoIGpiyYiinaonsL
KYVMhenLFcbD7kCwp06goAXhWDm4yx28WHP2sT2uidNQo84buA5UBRXZ//yD+ChJ
5cWmXATpfkNWXNTx5025+yPHEgN4gCd5r/XOv2TxQthSpl3Qxu7fqGlqLwVmTfxf
ty/hScc0r6vz1JIGsvN1yJZtFGAKPKuyzsD9+LLKrbh7VLecvECW6EH1sjO49GG1
eLnAKejx3BoL74eUwImcifFkRPwJEl+Vv9XI1Dc8tnxFztJidnzk2fVTbj3nUEz6
dUqJaiPb6Qo7VeiNaAXzS1BOd3+PncnINbwdowb2W0mkn9cQzaktkxzMOOtRurHM
PYKixSlpLtet/o2VhJnN5fheGJMC0dczhfaB96IL8rnX44ywPgNthl8edxH1+n1u
x0eheVzobH22KA3q1j7NwtS7w8CXQEG8tGQACGnyRaEGBxFLj7jpJA9zXe4cCZsr
Az9uk4reSQF9604Ctde5aQ==
`protect END_PROTECTED
