`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VmX091iKEO6eMoL9Uew6LnpcjPKyTRZvhnJj7f/nGO7CQ8TqYAYp5DnDKSEDCZUR
g0S5EA3Zq4fufOvSFALtyGssYJ+q+ctJLgc5G+p38EPZAKxkVDiLb/M4j4+2NSkd
+kSP+6+0jGOBF7oXYjNKfybs+Rq5wd/YK9Z1lBrnFRvI3q2kniR3tnDBjfxsAU9p
N9TuACQgPv4d0urVXBnFMwSY6Aq0lqmhbwQaAT07lCCVOMR6guF6V8f4guIOoNHQ
`protect END_PROTECTED
