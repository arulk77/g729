`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEA1tP4T99Fqy3softX0L3kjK1UCsT04MhZMjp0CDXlp
dRbb3fbZgrT62O8q5+MdWsR274UlBMVYK+hLC1/R9/Zi+rfzg9qCB7w88ZouY3aV
zmt/YCNTaJzEtlytN/uJiuPKMIhRlyMVqNuJDhH28S24pysVrbK+T+RK81K/4A40
0wWGGk7WU/F+Y1JYO+H6F9CEQIPMhe9BNO9vRRdjuStJLq9Q1bUvErTlrOxe6f5i
jOmDzKzb6G28mr5IBU+vOJ7Jufh3zdguSZaTODgV5EWLJg/zZgj6PU91DZwi7xdv
jTeMGWsIU0go3YS5PKfHmTDbwgdkgRgYSlNduxmOR8xc4uaZNMAojEMKP4dLK1Se
pc3CafG2pvixdQrKCiie5SRoBlmgO0/6clCbV1LryllOfFv8SB+9WW+MXfYcBLOa
wzKpWAuo+We3kY/IkfdEo+Dfl4hKQhSVVV3QIKIE24JB8NCnH35nZn7WkuElAxRk
NBwpmfOQIfjjQcu4iEPBjfwkavBzOoU1yCvc4qwEmRmDgKxNdxwc+kUxez1Yb7h6
`protect END_PROTECTED
