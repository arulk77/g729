`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC3dlbuLitKhcdqhzKym///kCRzWUbR3pDk/n6GUdr8l
0vQumHHI3r4mhqy8/erKbci14SKH5fklRRMGtx1HvflTXFbVqK9Jk1AXs3P6zVrK
zrPMK0dNwqMtR4EwCuvexZo4rL+jciJOLNfAhSjwQh4ZckUhFx1rr2L1DdH7NS1e
tKGjfVyQad+tp6fFTTUGQStiqA5skJv7nJMfYfDv1qBL2BtYUDVrmhbH3NngsA+X
/z2e12p2C5d4Qeg+pfzSB5PbwkI4YxsGiZBTUcEyK6e9DzSMJphEuS6YVlhsCYYA
GJSOr2b+YTb42Qowa5yt88AIOUa1KkVXEjdruqBajvD9x3kyMhFKTwpZ6os7aWIv
0uN9XYxFUrZ8WXR5w67dTQ==
`protect END_PROTECTED
