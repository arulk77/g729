`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF/vGec1PgEu5S0On62mm6b2nles4vjOC9DquNZCrQqa
DOqMBD9qZR5K01ZmLBIvd7iBDL4tVHmfi8OvLSGe/kCyDKhNJizjUQ6Kk9T9LY7v
SJuUFlA1MO9Y+mc8p82E8HoHb8gpujlInNP+i/xYhHiEVG9W8qsNo7TjeCkqIcQV
pyR5qSc6q8vGZXM5f3UG+6HgILv46/Lbgj5XGiIMLPnPX7qYqa7txvsZltor6dq+
MXMiIbswCQ1G4EtAl6kLY2dRelWjERyasoXg9HEUzkyoGW3m2EEG6WGg+ISSL4nL
BDUBLKaUyByCRjgiN29Svt09vSMQsqYKKeyvjpgZFqTw0+Ny6NTuRNQlO8lLXcPX
`protect END_PROTECTED
