`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePF/R0PCheWsqgTeC314UMZyDkCCyaWkJe8YRQMYttUx
CWoBPnxSQitycgm7kNIDvBF4dbRywitwUq7Al+OgaZ/tLhAaQLgOadr/FbY+2Kfy
8SV8Lp+k+vZU3b+ywlwqgfuilEvoyRcPUesc1tGHIMfRVzRCK3oMIzbUj2Brpb8Y
wqtT3rnehAvp48TgBzT79w==
`protect END_PROTECTED
