`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Sip/BA3IC8+uVMSPYSjbF6Q8xVFPeKW/V8LKdA139g2mHfDNm+QGLjdqcNqnngdv
SRY4ig1CMwKJVcQWGN3XliReQlJuIyIXhjoBT/djARdtPwO+25bkcKS1KQhUm+RL
xHWZ2v4wec6c/CeAjXSgdPY44Wky+0KCd4wVcc+FAvqybisax7za7ErWROM/gjYa
3DRLjUNmqZaS7eFebT4O/+Mkr1G3k78VkQaBbd8AdMq6Gok6XUVSEaDKGbl3r9hZ
nrB2E3Vmhsugu2YrjBx3oepWItqA52vpJEBDu0R+2mI=
`protect END_PROTECTED
