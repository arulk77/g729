`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM2gvISvE/iu1wquTwki5wZYRFDCZiqPJqsSbwa8w2Us
nEGs/2EKp064tHY8CyQbhLH5otiQ/LNDL8mv1TdSA2jilBlxzv4PgVJxySPWBqc7
PyolmLxvBdT7SpCIBv4j13Jk8WPuYEHh1Y2h6xYmuOUgIsEVD4BwMix+3ypZN4jL
/yXXKxgpQok3pnBqg6+dFfxd+RmdWvG8G+iN+YMOPbr61C+lGcdAT+SAuXCKlT6N
2L1dxWK9++yVLmIL9QHOnrSBe+O3xPBjUntfl2Wx6v9Wn6oN3kJmPrOEpLWdxzL3
85kcQNd2F4pyCoTKJcg7XWzgeAf8xR6g4CMNCTc/bNiQjDrcw2p1/RdbSshm/noH
77q89TgS56H++cVxoWHoiEQ7YZF7eCzO/9IiPDe3lzRWTFEdBKwDl9v2AtYzx2Vk
ULKxA+mdVSlGJmCVVO9OLM2cy1lkjBqJUffl/wD8W1Opb6sAyYDEPHixA7Z2bcPK
GtkCrNpZ/xKV+fRh7IcPGQF4avDmjAfUof5UA80gi9zZGn2coPwsiPEJb/lT6m/z
`protect END_PROTECTED
