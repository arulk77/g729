`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEQIx5e5Eqj7JDg0zJJajseZAuDeL9gbydfML8I8UKQD
VtAlj8tCexHJhnxx4zCZPr+xwgflpuNXVWj4KZ3fSqqK2rOYJIrlvJWgvACDPrJJ
CuVnOUVk8LPFYjW7IdeHDg3R8Ji5y3ZJlTKMUZ5eHKv+9xq53yv5sfL8v9d/gqPg
j5Wrf2LMrpFudjBGMGSZf3gv4DVFwrBtg4Pm/Gi04nwmDXVxTaxmcO/xEBbDLUfr
athqjzUhx6z4FZnjDp5ASJhyQ6YXe16OGiUbObHCLvQb9bVWO8xYoHburKYTZLdw
ve6bniWTntcy/pRkrEMViztT5ELFxGE91grjme23zROKU03fWthz/ke5bwWMHpY/
ZF1oJjmdJMpH4Aaku92gVZRipXJ0uCM2VA9amulYZLAbuplpKgQuR+VMDnb/3lNR
Qmxn19J6+X66kGmmfDhreokib9yBmf3KhZH/LOqAzyw/IFhCgl9/BeN19yAoPYYb
6sMI/7CRu00VDz86uKda/ccgjEgbN3b9eBvIb1iw4arxIOFUcA8ZID5R83fePUbB
`protect END_PROTECTED
