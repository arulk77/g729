`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveELdltX0Hduk7NfpVL7a5nifC2Qg9FPJB9aYBBNDxSJM
53fqaqzbpX8d0dFInQkGYhJFMujBGuqMZPQzz0Wt0t2LPnoLE49FPWyBThQaCYT3
RkgfbjT43AEIyl0odmqXjC5Q3pG5KUF4HXISvgQGiZU89WuCQI063vtLk4Q8zzNr
Pp8CEMc/w1tBBf+gsNJmRCAKWWsU5zRIqlDvbWYLKcp+eBHXtgT0253DO/JN838K
h6VJX+Sc63IKui6vgFODr5Yo7kBd+iTj/YJhCQ0APc9Ok1HwCzoAJ3z/3ve2iOr+
19nS98jRjvZ40oOhsXuMxw==
`protect END_PROTECTED
