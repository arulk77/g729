`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UvOW8ox1vtNTgOpbWXDkTofDwHhbJYilJBCZYxHvF4qxKgq0ONfIPzkkUjihCo9h
D+vDbWiN4Kyhcl+i170C+xBxrMgFATZKY/y/DpkpQJ8WmHoYDxpuFanUBMP4Prot
UeuEwKrVecCMtMT2Ned4j681zM8YTQABZ0tKB5dRAst31Qmv+VbgOlrU+qjUWfaJ
DUi4l+99i2yf/SWVoyv8vi+DpmLgPtN7jafHv7pwigTdStJyUvIRKdZkW29uFOXE
u/pzBLSZurICFSCYAGV2/UUEcWp9b/RkoOyJ/NauDN9OnB9/8SzkLmlM2N7hu3EP
3+bJtmLIHAt1QaLW60WCjlGduS2Bf2c4R+7OX/jhLDtMNR/dlq7EXolgXa+30v8R
HOcUL9zYjxcikSbdn9nhUmVUAADzL3kr2KYJznTBan2biG9f5YP3Hs+6BhVc/tP7
JMdkdzxvA0koSnkpzaKuDw==
`protect END_PROTECTED
