`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP6MD9/Xdn/AqBJY2kirWwnk2X9chGTgVb2e+Ux3fzge
finsDfo/FUkDBri57OE//kl0fykkEInysGJj5s4HIRUYx/ieSkJMyfdpI5Cy1pn9
NQGrrk0FErvXNkkRbeK5yzZ3Szbe+pkQhI+nDc7Ok91gTOSmEgcP640c68DIdwGO
vQq0Utr1NjB1So8aJC4snyX4J6Tzr35EO2lrcInS04U=
`protect END_PROTECTED
