`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xXX4VGZrw2rAKa6Dg3LzTq3Sd4uHh4lolzXD9HEizt6
5Nvk5z9nXw36dLuXOjgvTXEfhZECFg5ryNUnYBLET1D6tgLmFBVKdXfyzbiSL9kh
9M4bGDZxj0Ab3MBeJcBIJN+8OjolmJvR9g+MZn6wmwts2YWxYnZ4i2hXE+czUUtv
vIn8Pr5psM6zOyCBrb2NJeWo6erv6nj9M3GyES+/p2w54YT5B4UBQqI68/RZUqTg
qaRWLujzqmsPvmN9PDcGhG61gj4c9cfmD/kwtSEkeK0=
`protect END_PROTECTED
