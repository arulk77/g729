`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MQ7AUSEQ5OmQeM0sx2hitwtIEz+SysDczvXKS0MXpBhzBed3TOs2CZ19n0xxBot0
UjLKn5lWJGYsx3IDP6iMWRDywiHA1/MVsFbOzKb7/nEGDW4zQ1lgoiTGCaDGY743
1WZTQ2oBFwgBgT0TuwTB2w5CjJQoXR/mgQGnFkeHg1MzScsPT6IToKA6VlidosGD
`protect END_PROTECTED
