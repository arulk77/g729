`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGvIby7B0LExCXL2fUJ8ShCkjuIQVC9ndf+0P/WCC+qn
Ra3mWfEbCpT0xk65+W++UO8wKlXiIjxVBvEXxK7sHxXFJ3QzRDxNUnTU+SOYKTvy
0Lx4Y+/Fv/Mkt/gMSqd7T3J0FpVTAiVHYB4NX9MaDY/n81PEMfLMyghDgc+bWgJB
`protect END_PROTECTED
