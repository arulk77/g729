`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DzwGNjTtltPzj/PJO5VCQ9DXYJjjezLO26hAyUU3c6HEEofM9TWWRVS4SU4nc0mf
TXef+skXM4zGYAhmkCd85SgRFkoRL0rQnLYdOArRnt0ny7iRG556Ms287LAG+Cf5
QjHx2VmyoBeqeH4wZ/tdsJUsaKmIjutyD93/FSN8H0v/iRgzBQQxHA6RCWu3/OXg
cOXymwCRPI4S7VKwyF81+VPUUa8/oHJPcDRc8wIP1//240fR77FH6QbV2wfDfTcp
75i4lCwfQgv1t7cOUxXcdBxZUD2CK/SxyEh0KhnkxGIP8ELPymVNfBnBPHg+q1uW
ON4D1YWf7wxrHfXmhGwnH8oxiAPFHAZT16dgsxHy8k8=
`protect END_PROTECTED
