`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZZnh8bxlyuiSQrVnvuwKH5+1fT+UN8gVXYoIUDOlD1Y
SU5Hh0oi+yP8Ou1rcUlfgvZoivzeDT6o4lQ5LYI/x8NvXBUOHuoPPih32Xd6ONwA
0x0ktQsiRL/D6XCrke/WPFC2NuzTfgt6mM6uNuKuL+yJcvlpK//5xBWVyQVdvqtl
PyVv7kfidkxp8OPsDRyqbo3aAy3ZtFW6ITpZ8X+IcwXyV3nZFU+CP5vSN8yuGAQy
esTfsHVlDsOqQZrO1TMurInHoHXJeKYYuq4HklpTp0pqYsrqwt6epxlu3tcrJjvf
TnTRpOX1lWjFrLKpB80DWzI6siUXAxYjnHLT0GVA3IBfc1hYC/aWIeTdZN6LPIK0
NeOofgUQ9p9s7nhPpFhxQJZCovgMMH+uX1693O0/RmjphOjX137rdIrGztkgd08q
i9gLjmXpYWHfEG+jbpnM9OsPQf9dk/hXMDjn5Zi34oY1qBisYWmgK5SuakVPg+pl
PTrE76awhZjeXJuQ6IxqpO1uIcYyM5gTI+c0cyFJ6H969Ca8o4I6wPJYkmaszqVn
puEhzK1MZuR/eEHjJdaUEwngJ4MFRwp9y3BnqloGC7u+1ariohilfV7jOSnkiLYP
YkWyOo1fklUDdbeDuCo9Sn7QHQs/4PFdB47mVI6nRvEehQApiUHKHgMIUNfBQ2Sl
wMvGXVsKVgNlbBQpuncNZywdvxJS5pKNSYK6LPqh981wvir+VoQ5yeUr7yJrJj5D
AmKB7y5i5vmdBxhITRivhQ==
`protect END_PROTECTED
