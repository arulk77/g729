`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SrAwW1qQJKBTiknXGU1JXJtBjOEjv17icNGTn7snYDfhSuYYrfI0jZ4VciCM8+r2
uD4o1wYYzYaHoQe/15FWlUbaUdwL57rBuG059Oyqe4vsz+8zRhyPZghlvlxL8vGc
iATtyppPW/BFmoXUKtmj8gEENrH0bCIzBjVfpdhkasVypRk5UcdNc0Wix/7gvXDM
qYQOxZ+RDliEgqjeSCvuYlmJbgkavgR3FDbLUxltXeU5o7HBB5R76jx04OB4dmlm
r7M7DthOZmGizQhy/Nl6+k1loP7AH4wAHmCbM+gu9oInLgSXEEkwWKO2nNtAR9BU
nZnqyeblsiuXvd9qn7oaONFZ1lr6q4aeTrPO/0FpD+4=
`protect END_PROTECTED
