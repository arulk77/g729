`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QsIdsVJhb4CckeOxRA6x2dQ7bBUibcKwKdZdeeFjE8F6pCXxi+Y7loFBKGTuDeAz
apwBmX6RidgGU9Wl2LpR+PU80SUYOErc9sEpOM7ATJngX7WfrYEJ4QTXQw9SMmhz
sI+kccHSEytmXcryTEQ7iiOUe5HNoCk+o5YSwyzbs35un5ycOAYIIgTk3LrHPjvK
SytYeAL8G+NNWvdmxVAA/Oe092HSGoASEdOf9OPUFXYcNIBz4gpuoSvkfFgypQVv
8HqPHXIMZvcT89QIJLAfSGiYj/X8x+IX0DNfLm7QEwUvd3timCPbLL+6XJd50a8S
vMjpGf0BU6oKtEpLFO/d5nfFERyRP6xTjordJqrXbjv95XfCg/AWKz9GLYsn3svw
Mtk6KOcZEH2e0HnWtaFF9vdb8Aq+bhobaEQ+mt3NU66dEEbkb5OSXyrUif/gwyUq
bkO6KXHKsSrPrQIeve5eEw0C795oE3jwieVMNdhsAeXEaV2gGGJEZwz+S1o2AIWI
NlLGpMDcf8XFPjOWbFkmNAnMEtvUwa+ZWHNzAnjaX6HWeE0L5QilWXJyI69gBqPQ
GEwT7VSjsPBzEd/1AZ/thRnDttWuyfD5Pq14JCndWTjBprAHOmOYs6k8nJAtSXv0
DAsIgVbbHuKWJVGFeGVkUMw7VHaERCZOPlCoFwRYDDhXNJCN5ELCw3hboT0J0Afl
LkQk2YdOY7DvxmLxpR2pqX9X9SYNAC8XT3NQ0Uq5D1DOeLQtJ08+H8CNVGdAQW2s
d7gTLHA+DcJLiLlDKGfbv96jWoc4d/UafzBuJMw5eJ9KuE3ULgQBdMpOBYz0NfnA
Ys9n956T+Or90PUr8VDfnFaRVcdE3qYzzqh8EALWhwQSblCQWEFkNTmkVf8vsS5U
`protect END_PROTECTED
