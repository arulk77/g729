`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNTAt+gE+IhNAFX8lKgTvGqGkcdWVG9oEAR5p35iYRGa
vllYPvbvp+z5BP6zuPKncMt0/GenGAuLrUQeF0gyg1rPVU67dzJ8cakH/i1QNrVs
Guv/gTyR+BFtnyFues4Tjz5lZpQgGeYwjU25g7u3kQTKumFyoCV9eHikvCHkYnrF
ec09KdJCrheBqp9QEj14WQ==
`protect END_PROTECTED
