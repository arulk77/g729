`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKtM1f2mHzS8pgxje4jMXwE1BkxU/Wd7eyaPXdKelypw
JP0WZkq9moGCrXEkePF24NQhmFwQHcUS70HvijiYGBUFm9XSmvrRW0fCzACvfOq6
jD3trpJJ9NcxoMukfOUlZQH4T/bM+l8+JK2m/jUS6GKdQ/A6FpO9ulmclDQBVf+2
IfSOLEZJh+4hSN+Vz0sw8olF08anWRmJ/pn7sQsEcXyVC5Zk02OVwLLqS0GGzGE8
PQqzrpupRIxnU6YzQMAhKVKDrp2z5U0A32pgly8jn/u+l8Y7Keqo/68WC3l0xrg1
iL1K86+XzPid6DamE2pPyqMyTOiSQfId/eMOoQBifgYQipuhkQcjBo5qr0SS2WVy
6WP8YLHkDJRvFwDyJFiyPmytJapbNlWFHevBCVtfESgHXdFtkDBhgQoMPajKYHHQ
6aVYLuiI1kGUQbIlA8kNFdWA3GiyHp+Cgez+Pmtyus9KCz8FMVGeNM7Bm8foj7kg
ZB/FAA7yYBtJUtXmMM4B89QijNMIXWdNUQV7UFHlk3KCsBGkISBmNrFC35+bKZRO
RI+N2jmFD6uwPgVxoRFoDiPhS3fjWLPvUypQOCiQK/Mr0KzG6+F6u7HLliqBStFC
wwz+ARDujZABFr0FUotmRougb7Vu6u9kmmtqA7y/l7f/ZXafVMK1t3+F2ASUgkQw
`protect END_PROTECTED
