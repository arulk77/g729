`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu470rAMRg3cv1G0ZJW9bLPh19DTMQLnaBckkTTJR3hyJt
bovokxAyDcNZ1MVr85QrpP1CYKH5ryh4lVtexhUY/cg2+MqhjEBPFhnaHjb1W8av
g595eQHAnFMpfr8OdzDVnn06e+OO3De+gH7WzYGMgareysM730mtHgS4A834kiJY
TJ66LrAiuOnOLAkYqxwh6z3SQSLgXrevqFVQR/fDtoQjsNoce2JQK40Kwo3lPS/Z
RtQLPUZe1Uzd7zj16TH58w2mWNDAKjFT64y7yXanOAA=
`protect END_PROTECTED
