`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePBIWWZ+sbtsaLxhc9yYiGBEsFXNwRgBin19W155B4TI
mrpsztHgwhs/YaqIHVFEOdzGf1Oa9WZl/xByRHjscejzVjItXwaDvRYQHFbDyBRy
6UO9i1OwePuNrqQ4p7KwtodYC9ilXEg3trykhX4eZaKAXgoghKM5lvViX8SFskUg
2boPWGigHznHoxhf2ddZdb1EEHBpwpwY/arCy+ohTcQaQ2heQKRpJNmRosiDJ1wv
/jujfBmvpI9i4iTXUh8edV1+KDIfTPD0ZU2MDZgxGxA1N/Zve9pWSSwl58CHcum7
dLwcb3nKhOdCsrwwRP7i8YBcI/4VOVLsfNWRWgmFo8u1PBDdcd0ySOE+62+MphII
ggc5PlTKrpYekvW+TLb6etbs/QC0IPLiAu0jRmd8n+7hDcfhqtRdJwypFl6qd+5M
T92LUmF8thqpTyNQhsA4robtjskLRZHSOgVyvyogEESpdGf6oWlBl8oD6k91K0WQ
WlTvL8U/M9BQ/9gGkquO/LJllpklw3AnGQvZ3/0ysGx6aw5UNL8c+wVnpOAZTr9D
`protect END_PROTECTED
