`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFtKCt4vwLBys0bf+8nCOBoHwPCMY4UJ6VbGjhdlKXjt
+sWXgdUwYD79qsHdN27TKD0iWlWudQF7g+U+nweA+iXNL+p7jKXm5WNdUIGQvsPx
fHLWKBZOGQuD+1JvUmDWHc8hw/y+5cPLSM8PXhORhI5aTYeJSJOqTmbv4y8Gi1qO
52fd5yOQMMGHMiHyMCWAsVmp7vwjGwpoUCBT+KUl0gSa5kvig3bj8s474YCx9bWz
p7R8cDTmZ2qOynASxnc8OZ9yu2fs1kAE1TqtskeGxKvpSEMIspszA8caVlTf5U/5
LkhIZjJJ3fZYRsnQGxHCgKXeF+wI8keE1cwr5alAMK/PPf4UwVqJ4rUxf8w3nA+3
fWZZYe/+yLu1DdH2gjg+KyxByDqUelhiJE+D2iVCtuymzRvBW72yQYV0k12ADQa0
YWA3uEuqGi//2hV5NaUPplBMiF08x4ptPH9/vAqY+a68AcacxUSlv3azqmGXfboJ
FYJKO3OfukeZpyTLyAZS3oeD0h4izef9US3ViVL8qyTGY4tCFVz+OkU0Z4oZOWP9
184rH4kGNcFvelXTgOst4i574fO13ptSyJ2Mw9ypB/alkpwtt0+aEeeQRnq237M5
`protect END_PROTECTED
