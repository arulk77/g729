`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBP1xDTHr8YPmZVl7so5UUTRbGqaKSOoyNEn9ObWVN4L
nLhUoURjdJf8v2lJzS+DXK5EnzpPpP8lRnyPDKlkWxJ5sC17PItS9ElkfBtwYl3i
LSv0wrDG+gIS8hfQZgQZk+tQ6eWfBENZalpgPt13Ilq5V+R4pOQXphFQMFLkfGMM
d1pjUXtd1kOFNAkDa3FbiT5dHrUrH1SvJrAoiEq4X1F0zSnstpjLcPjy9UBkRXLQ
l9I1MzUquOFNEvpsauATavptwtSPnepU7DaqYz6Gy0CN2NQRVqSK43TQRYb/u5IY
DafHsMHhYHxyskgHhPo/+cgzB+2EpMOxBYwcESX+/3rn5aaIbAzDcH6b3d4IYRIU
RreTx3IvZ+kUf+oM5FAEeaHumIhT0ZgCoboegWMRzwn8KgphIoiT3HDbXHln+j/Y
qYi2lX9+dlYLrC7r+magDxajbu89VR3j6zS7v9dp09ywUoGz0mA8iS5a4H7nUu87
qip7sIDXRnjoA9nXSL2opGVCoaFTW8TyOBaL+7MHVfNumGvIb6/2a2KNeIN6RieC
`protect END_PROTECTED
