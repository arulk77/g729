`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43UtqWYMcp96kzCZxdjPtS/BBEP4iJa3AzbQeNKekpfh
4MpFjjhLtXqrUf3dOawt9krvRFZtjKwCKEm0bkPcECqFVFmklzGRotjH6U/b+nFt
kFBPgPOgndlDz7pIxH8MckCiKvIWYXl6/f3ECH5f/RttjQLQXowlGEB8itn5gyYX
kQJ4M8m8YgCjTc6miZdpcxAGA1IZ8yAS00/+tMmY445T8pI43yS3hGc60sS0zXF+
OVM7gzO8SwE7gTAgDUDnslRn+nmGVDfoleWDd28BYHFrazvXRoEqjNYiJ+BlJMgZ
LGUpOlQgms6YUeQyjwIsyaZcZCt8wVeLtSDkbi8GIAPZprjJsXtW3WSSpUHpTx0b
ir6RKpx2FKSgC6BVbPASGA==
`protect END_PROTECTED
