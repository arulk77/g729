`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDlRavDx0EkRHnf6hilctV82tQcfWWQcsEaeEDNs5Jkf
R69g0jWVTPqbJ9UE7NPeHB/Pp8Wpf2vCRiC8nvN0MP24y+ebdRvrXdxy5+r75WiA
expO4LSFwLLmmI8laGg3t1yRXTX52EOIfl95nRqtShqpcwLtsl17eZvMW9s5NMLY
VHHFZU5DCOAanYs43DehwYHadLHekUagcRQQh59L8KvPiS6ffk3KbAKW4S5wCMlC
VBPs/MRUhSZOdcj9y5hqh3Xqz3j46KQvtXvALl6WRHppUluwcwFLpFWsIEE5XBdB
0PcqaGnSOyVIg48oVZloXKjJApMKYk3aaPBTKYGirnkwSOijBF1CB3Xo5XBgkCos
FCdaw/YHedYaZa1RTSIB2iqKhJk7CMzXVtTvK67/TfFcwUH77hhqCxK7CECfVnye
zJiyvQyBIYPoX4MqS4dV+g==
`protect END_PROTECTED
