`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aX6YOkW6KG6TGB+WZXDCJ+UwmfKaOtzb3P8EHbgVKvbQ
wiAwZ/pGDZJW4WF7sZn/CTlAAF4Nyc1fXc26O5ChcWmYx/edC3Dlvn8umBDXUvDH
hjcllWHv4LvHqW1RIOSvHNLq7mk6E9Pk2f+RcbYMF9hUuNDBrWDb44/r+/XPCKX7
Hzuh8TciFIumzM3QsAJA+LHZpR0xNiOK6nsdiLotDdGAE3ponSN5Tfq7DOVrZHy6
PF+LL3rXZU9+kSzS9tzF9FsGp8x9F2B8FbKW0NRA8XQ7dhVzmbddYxCPG5/9Z0MO
A3ZgX1I1+0tUzaImmBalgdSlGTPf7h7veSlCaVtHu6ElmFgmERVS+H4SUHkCa0z4
8HJqFyXIAXksTyvwot6vh0JpH9/OAbx6pF063vln4Ocydb4dX5AdLX5/iOPSht+r
gAyRkozJ9fOv9wICfr5EGsmBogAaPckRLJD3zm01ZXqmhq0VV19ShlklIM1rG/8P
4jIgUyqzPNYGmQm7I0UcuTjH2GXvKY0GJ6/nyNAth58tnDhRwfbOSMDxCyQ+nk2l
FIOMamULrn2CWGFw3kkEqaRtez6zfLw6eCRi3ZiLcNfYXyOa2rbFujdXaAS0PLFQ
LiGNHQpbv7dIIaDIlho7aYKLAt5QkC9FKazXMgdkFpsE4uruAef5sNHNHGZR0t42
XiUtUbBSuaeP0dI/s+n0utyUjO/TZ/UVKN7RL6yUFc3LgiiswHhehhV6uxsI9cER
UaEN3Zhy/BzmJCallWme6WWQGl9CE+/2bFzY2BAVaSSxbrm4pbc8+eizYQuUPLLV
hNlO1L+uXdZi0ly4WnSVI8DyXgHvZerjfaM4eSS4Bq5nOzxm/mC4OgBnOMeDJYyU
X8vzxu5qWJunBvR4MXtmprslbeGzGK3mrIf4LtwttEAUvWgY9Lc7Mlj6kn9p4Wig
ymIkkXteBJwgfdHHksnCbngnmsHTPAGHEQAfXiF4CuvQr0rMrUcbqNXm93euWztF
MOnypz2kD+bL2Du9p8eXEo6Tf1cucfOVwbZbqSjfUGP2eQfDoWYBoCv1hFzjEVnj
tZxRv42FY08kFgX/TmLVME8KM1ufokIPRVhm6BDJrH9cVPMLFU+rQAsTmkA+dxaA
maPhr3MIk2B8NiJGsmPAn5EwASM3UVoTUpXGw27XuR6O86Yg5BJvGckekoO8Fq0o
tQDPtoqo1D5hrX9GoPiBzq9x5wx0D2wqUPZBZRgdWfTxZhLywLvqXbHydYR47H3q
9TH51wf3zj70+BQErx7CjI38dDi2B5jx7CD9PU9KcGAPkgJ5ZUFwFctnl2QXbwoV
+En7OpyseM5bMd/kl9I9HWhTANsCs/peyNZDx6FEagxlAdg6lHeF6ZXwypPUrobr
cs0AkhRk+Q7elXJ6c1B1eJyd48rO4k8VLNJGSpDjOnhxgDzB/3lt6wll2LsKT8tu
tBGjpq4nx1rgpGtAzpNtv/UKvpP0h2JcIZBOl6lzA/s17wAI0DZsMGNpiskEWkGp
sSBJ7nNjTFxXPHvaYlDBQpeCtYP1QfhltV3lo2r7tnxC/lfYRNKipY3ADnKOX4XE
BaKq8DL2RT4b2ZgdYhM3OKwF46ZFNVpQUWy+H/EGsmlbOO2JUGsh5yQWMUw4LDIO
WPtjDZ/BFuB9BOrpaQV0kTadsFv1Dfs+CY1xPAYzbS6F9oWMSFfOeHPqzZTaH8fV
upXrWUxshgySx6xIF6FvIuFXSNbnhHxQi5b5Ruy/3J2k32a/prL+kCzAf8taCqF2
DilYSofBIm59nSbGQscGI2bkpGL8yR9hgt3t0VUROOZlwd/6B3vYV6V4I/K9jQch
f7pG/MLmhPfWOSH1XcbtEcbkKEqy05WNsUQiOc3PTddi4fen6Zr5HHjMUlGnvIDf
EJdY5jJmw46nJhZfrc82/yVxDFVBESwXvp/EKEMRKpEA8PrpKbg9k43CXGokOJ5Z
uYuaPyy6rtjBEYxrNOi8XBKMg21kGjPwMCn6n+PqZtjTPz/ypxOxO2dnosj+L4SA
VZbos0eLEhlgOZTWHfRTDubryZG7nPCYbb/ve/6mSqh9Vfc/VdtqFRplEYKygfxR
97S3/BxcGwJ9FUkzMBHaR47Jmh+ne9OKr+i6MAGn17XksBUgkChTk7krnSNQeptd
CC0C0/ZfDwZyPUw/7vPHqAPnPSip8a30DrAO0lRa6J879UrEhgoQSVvsA8+nnTbS
BVIalmbyaZrGxNaKfOwxnKO79te+Ad3Nghjn5IsemT+Q+h899YCbBF03VGUPQvnx
No9GqlYqYen/3g648wFP652+yCYIm7KSq2vhvs6mAK7nw7a580vNtrwgwOun/tOF
KBkRq5A2ZncAkdSjJg3PK0mVDdJv+E0lbofgig1NRUXHUhMKPNel1eOnZyKrEvgP
2wP3Ni+gRBf6hG9HtB0H0znzLA379Eohe13+IrJYPh00fmrWX0xjbO2GAbWhy9Ji
YRpWWSZozhnm2SHRxpZDZeldD/FJh73vePRckNlv4gCP14p3nzQCXq7A0T798hJf
esEynR6oaHlxq06M97sNxJsgbMLEeMx+PM5EeVWIUJyj4f4/E3r45qkpHMvMetKY
R02C7xpLOmBcODlpLxpyhqWx1safWhOPuCiiB054IfdUwVIXgNgv2ss9WqNpJ9oe
dDwRYyG6RBUKhXssMz8epwbIKVoLP28k1a/CZe2EGOpa27iFXJHDQDiGS1PGGIOS
mPrv4BdFdLqykO+GMbTtCeBoAjCTs5wMXB73QbtMEjQeAZg4UxDc4CfeH2H9iTeT
I3j5vxFfHmabhwgfdFfSx5KAhIfxC4MAP6cld06HpPY/pU6cFrUa5a6ZZ+eBcf1N
rb2iLQMqtdWd5AgvdOtFfADcf5otbPsUGFymLkvSeZ+Z1eY4OvmD4kxXTgPQYLZ8
NRujEHBlYBGtKD4uvJmmozaxIuLoR0As+3baNF6eqSDqnlaN1Lftf2CRIJt1bO6V
VbWzC/YmxcPs1m2FSLmM8tEtLI8SRLhWZed1pLKxspM2CQTmtzZ+rPmWFFU5QVqp
oBD+w6Sn9yW2JRrnRmA0wnUP7sfNOaK11oAEVuR17llhYRdLoEYP6Wp84skkEGU+
B/HG/wFFyUrSrl4WQ/cYWmaZRXpfGjp4e1Z/c6Nc5/zvidd2KG3Y3tSziE2mQoEy
fWPTX8pEPKpzo3GhnRVhk3rOrk6PWrVovsEQBlIVh54lfxBdENZ5yfEk3iikzA3T
Ji0kJUBqgOUO9781H5EVkflvb5e155qpqQQDnjp5c8eKm1QWR2vlXOi5VxSiB/R7
K1U93knmv2UxJB+u32StdfIHzrwVz727MleSceiJ/M1izuGnAP4lazHO69gbuSJD
jTO0nC16ch/3zSHrnTPN+NyUznfCwSEw93sjydBsoy0SD14bqwfVVL0els985Xzn
pWz6O+vNeheYe3hoUafQ0SQ1BwPnyUPtCeQAyCCHf41sbxIVuu+o+a4mExJg9oGD
H0VflVNB2h3zPGqDv+ISP3iFi3zpU/pNzPsurk5MJwtZhsxV25NbF3IOb/58o9R5
a9sSEFU/QWJPJB1Mdw42Xyl74V75xiGlGAyE6jS1vH1vxA9OQZoZ/KZJ9YQhBSeK
TNi3iE4SSy8Xh98DkE51XRj3lwUcjV9DL26iIcDhmjEs/I6Re1BHkVFPW8KGumx4
x89ZVBxcy5OOFbdE4jq3V22a7imT4XRvoTfVKP9b3S+H4IWXNDDTq1Z2EPJvm7bw
uaeZQLg3z2lHaKloZIxG8bV2wS/xCieICRHL/RJ4/nV6mbzN4EGRnis4MUU4YZIJ
Fu1IbFMbg3NB4GfNLrvhvnR+7n2HP50Lhlu7pAPWOUp0EX8prK5M+12zyr/UX6YE
/XAwIBp3BllelKRKCFF9qeucnnXE5zKJ+hQTJWP6sJB9E2yeh6uY3Sk9eOwxNm1d
v6EjjWtXLnl2utA6qnt+ETTP90nmaSupnnjIwZCwjgUUo2URSz14eTzGKsk8CYim
fMgzaVfeH102Aav+wL6Mlk+B9VGInD5+GvQK70eTYw+DIYieqjngCgXUktlHpGmv
Q2NkGGoqcgJqR7V+4MmkHEB3Chi60FqXi59m0WWhFJmyGtGo7kqvoPB1Iz1Z81/S
e0Z7XwoE3fuYmKyeu+sf1mPzmaKHosCjnd8I3ngGjLMGlJU9vImTjplmeRi3Ox9f
HMJehV3desMGZGqOU7HOw9n9mImjZqrAxn5343c3J5h3wCsPLBqRK9FWj0Q+sCWx
wEiF5tG9mKrcbbg5zjOVn+fRUZ7F1xjjIxAQphakqEQ9+xaTn/6niY6bJnBpwtb7
nJu2lXBKwNg/hP7LDEQAGI2SMQE0NVd+aqBrZUyoG4OeZ1q3kujy+0lb6iHYidpM
2hi4asz4O+fEdYJCnAbxqAhSmEl5DUNYlf/AiyYv+xKGvOcAbFtLNVYctovtY6lw
fugiwRe9YG62zjT+MFnSSsbrfq+apsCys53SBsOuzkRTUEpBOjFR6JNzIM7XiVDc
oQkqE8PKKyYksNbqXwoDTH/7WcLJ81V4k2NaLGdr29iZs8VUgYrd+u2bF/Q1Mg1P
Yz0Pn6RYwlgOYeC1mlc8Jwf+cxI/TmKtpKZdXsa5c09yKNIZCDEoxvvgDaDQtsj/
NGadxHpIKVNBscISvyqhp3/b0zNEamxtraoExdf28VrVZJ+EpzcZYMPQqJzyLIO5
OR6rV9rlCd/rx+93IX8cUDKVbTmyS+FvonLSgvjDPqDDZeODXAG974G7olIIJfq0
RZw7y2ey4330XHp3bpe0YickeW6uOOSgDO9JugzqogXzEurTW1WPi+tulRzuSoih
C/kPzmo1mDZcGRaBHM/l6UBIO2xZvVRpq2C4ilerCgbT20bODPh5ySkwvxNqhp7B
WVMD3p6bgr3TedXp85XtFVZfOES6NPhF+KKSBcs7NpOjtnxzZJSzDqMkGjQCiDml
aD6Obsgddnu1gaRsY+C6rpptQzGpXSkNP9mUAEnWCccOeNAp0sGswP1/M1yXP6tr
zf09TiSFZpnIad81hubqN7Hx0oe2uPkVN3DqLrw1o39+8/C4BK5SAijxUTEeADvl
iIHPdFfsI+YOgjOsvhOCQkvXmRplOM3pyzzjL4GC+w8vKqQImAU3y6eWWXOofOYE
ycoo3/uEEZXqcxKc7nvm4wNRCauYqWMegl3RQY3OwrIaR9A5ZxZmZU1aZNm/lMWZ
TzfIuahv7Sg2smgKNaK5udipiwVShnx9pCPgUy0CMc5oY4ejjl1TiR/oyzoP/5sN
FXSpyEUyfbW4uyozMwDrCzYpXcwmmuV8J1L5Z8YLz1VxlFvKLy3B7eNX9gebLqPy
T8+S4cTWlvDuA0vWHekknQ5m4ZzcaDIZ0hNptuVyUceA4UuRoYISYPBZMlmPHWEv
ZBsyRmDEC8QD3CrAUy7Q58dDP0Jz4FfxH8PHI23Klx6247d0w2q63ZrsZWABmQ6P
SylIKW6wuVIK2JuR7OCSii/4wNVpdwmA0R/SiraaG+fv8mKXtUe1+G/r+GJDVXyp
4GuIAgS8GBb3otSg4jy0fHw1WSlS+LRlaZv63bjXwyubnEH/dBU+Zj01LRbmOcET
jU+glywTzj7TTFRNWANqDUaNJNBvrBpBKhqv1QpIdL6kVeiguFjhgUnLBIUG7iGS
MfS9gYzVw/AsgvnaRh4+PEORxyFOabvH6n7m74nPriuyX8dsoLG93F4rEIwoajvr
VjGgQ63oVg2Oe+/bYJILd44UCXFixRXluIX0JDk6AlyNhwuqKfckK1z3sLj4/Chm
qDtpeiHCEgheVP8by/i7WPKTZfyU82E6HMxV4KUkpU6ddVh4v1BVwclLuMnc2RZd
bmIt2sg5lIdMZz55AqKF0toZenyC6JhK/b9Ld/e1yxemPaRIxa/ExcITTuwhsP4Y
aQ0tayMXgldCqiHuQkACpcpvO2toTixw8LziJjsn0d1uPkXgcen6A7WXway+cfAO
mhCwY1LIu5FXD8oggEjosbEnKIoirQM/s32p7RCv6aDoiH7V5n28z9pmm2jjfdhE
2hpe/m1lYd/GsZya0X1aWUtJPOgU5glHGbteDW7HqUcImMfHoPjz1WWKGNM/9lDl
T/VwPWERCotLvhtRG9vTSv4lnCmalaiBZbUFpn6zya61l0ZQD4Afjq+HJw2UChQw
7w8DET5vQUvXNl9ArnFMfZZk4xw3y45pLxinqjdNnPbNibxdjyZXIfkoA9ib8OEJ
olEzse/I+NZHgRVO0WGel1wy7FEXAROcOebyI6k06clcKDkeJ1tYUVOahCcFY1U9
6DlpqfH05htZQkWjulkCwHdY36bmCG4ht7ijR988y+FQlmT/hvuW2A+cUGsPl/UG
CDyLB9YrMjEQCBGESaUU9+BNRWnhMCXpqo4xwrv30vykPcF7le6H6zPya2cWL+eW
xN66qnKHNL4t4ZEVzCEi1qjDL/ZPt+Y5gatCdiii8oUpMeXfSMEwMrA50KRfFoaw
GDyiszM2ArQZQkdraER6y2BCD+WkTg7bpHu06fvi/XaX9w/7/4HLdRBf2ecI8ahO
/HLNlRxwklP6hpUCJ3COwdDBYW1fvVH5cKYhc0peaMN0NnDbVn8i3bIpB13hxi0J
qy1R7FCK9YgMmbXDyt6jGyW8MVpfJdx3rSbuNjE8KX6vIXyQh+edtp4/+tQUNgKB
9LAz14syxIbAmQYdv/7j72pw5dX+l0TqaQ59BIOs+9fZotlNHAOFSGNnWG/MJ7DP
YtuADx4nuZdb3BHc2cfUooDG4piiQOVvfJpsWCNMj5SzitXTjrptfrXrdK9/Re8b
d38oImtFJvedRiXR5+TUf50F2XvB3F2sArScrIMHtg/3iDWQLCZtcK8u2gSm27WD
ktO+2At/PVcA00kTUMXfHF3UIEbdgeUIVcWwgW7ATrQPNcaOOztQfdz9MXIrbRol
d4St5HcdZzssD+zYHlvg+RgrLGPTJSS9GxOdp2BDzKtgVOX2VpFN6JoA/H9/fp0h
vVAxhewtvFi7kf3LJ66Y+R5YULJ2BGoL++c0RiVeqY+lE04eGW8cPgb+XjLhedAo
vU6zFROBAW0w7P+GbcDJE6kVTYyK4s5H6ivcQPqNRfyidrGna/Cul+sOhpio7zCe
IbDZ8v/oLO+Lncttzz9kIbIkjuvpWlsvAb8wsAQEpucsQjTzuCF9LzDE3R8s9q1X
86zxXBhJqFTFNb8zUIAbBVjtWh/MK9raIA/O16snQf+aWekrhntDKgk5FTHewL+i
2IE8/Uf0HhGBFSYyCXOjqesu+jz0YniH5w4+pUCbkkJ6nl+Dwva0ZefU4JiyhSrX
O3YiFOhF+3kyA+w+l3z0VOLyhisF0zcKw5aDBDZYNShfukmtkj6EahhaaoI4wM4a
dnTKk9vC6UJv3BDJ+P3tx9JLr8XOR33W9S/MOR4Q5AG4ulFuK54ywBO60PB9j/aH
lvpnfVmQuKmMnBlI7rfzvD+Eso9hGMVGSlq2oEa/EYuLNjt3/MNjCQ2W6XqPanUY
pZsoG+fpo3k+RpM5Xk6O1hUKs35SQ2ZFBbetJ1pegI4LojB3PKlAMGRYDa/JLmjb
oQiZ6mIg161P42y+vjfI7Y93BDkFPpFXJ5kkrhVAfjcS5yrO5Z+xD9Nj3qXU8tl6
/1X4H/AKEQ9XA4mOHeSSyQJ4KEU5Eb/WRwTYvA3GxDBll6ga2CfVgNYJ2CAlhxxw
SGJCtzVuMdHNQIqr/5PcwdY9d59JFH4d2+mScsl3zJalIROj9mjjTzPeSYhMGwlG
S++726pULasFT+QXEvWVhCmrhgHB0zXZaRXS29D8Z6Zm6AMwN1EZtxZgFWX7l7sF
JrR6RPv4YaY3IaefM2ZuxtDxrYTO5KvLGesosN437Dadt3jqpP4hT4GQ4EnFgCW5
eP7F13g3c8WSD5Yz+S9FCepebNZJ0oJPf4VVkSUOjn0CoijxaoAVs/nwa0eYEnPX
0pCw4fHdjmvgfXKoTQk5rXwG5wA69j0G/XsTLj1ChuEV8MVBLEHyzGAjdUY1Hmlj
wUlKKQhA1rxUc5sktA1/TiJRPvhf5Ia8O6MAEYpGduCcbLzVm6XSbP+gjxm9LNA+
GP00+OpwGic1SCyUDZz78Uj4vCsxQt0S1ujri2fcif6n3sMgPlF4NdeMriWJ6QiW
TzC8uNhqoilqYmVARFpL4M1sljfgtFwYPHZlCxNlAv+sN4cBnvqMYxKLL0lrxhNh
+j4GNH4wT2ulLZ3UPVPNgCW4aGetobx5hMmPoL9GN41Yn1vvFFcyASylh+KPeJrY
VmjJKvrN1sxzjFdpi+/C/3uaSKtPwHY4M++1SE1rAK1FgNRvwZ3+6WWvnokTWKmy
YR78pNRaDIsfLTtmP8/gCL9lKHJZTUbLPS7OyRCq8bXDdjxrkBwF1HEVG3fU7mVx
xeEhCK3j2XQ04BCcWSscTsNl4XIrdrU2iRi/qb4qjLUyFJx92EiHoOMDsEwJHi2E
jAsskXp6iUKHhqrweUTkxtplQj/tjMCwkYVx5WQBObpqll2eiJwReIEcAHOkdIbC
XdkSVhXP0RBuNcMaKAchxEeSxtzJApf1O/8XNmcz6s74iegrAjIk2FkkcLQtUygk
3yEtXyTfrMW5qTHijM4+UJc8qlIDHlb9TqzAtOL2af6s6OXGEPKGP9IKrhduWGPw
PxH/7i+Y9KjS+pREL8GU0k/FqH0mRnvuMCkmJP7sxOw4bnY1ppDK+TTiIVtwJwJ+
ZQTDQaJBiBz5tg+fMQMF2ffzTfKXwyO2MMpXk93+mRbVn0S51mKsD7+OGfFT+U4F
hCRVRPNK/Ot+Vzx6kEkmUxlggGIdpfSoRNO/V2nHGWCk9ynt+EI+Qw2MvCXOgl7+
graNILHpR8Qo1o3itWEDvVOGOMBe55bOkpVMzzUCQ/GzEN78hKmv9SWZ/FSsocDy
6dqZDzgP/vFRWTTMTUXKLfatC8wsxHwLA6W5GAsnjj2GZMbLGN6Lc1cVRiz9GoJ4
7fKiSasDBxaKcyvkLHT01/4XKHdrEKgHgyRGg+sA5MEgOOt7zOEMDcauP2VtJghT
tyMJS+3K7wiv8KcQeOsquzVjp58emdrvmdu4l2tG9g6KabuDI2H6A5JMw50w7mS1
XvWt+yZJfpBd9wtHs7gDFg8kuKPhHAb3lJuZclEx+cmnkcPl1kcOWUC3Rg+K1Dp6
+4ilZyrR3UAgRmqQDc5JlwRH1h6GZQn0TzX3mdv2uS6KXKI7VZdruPqL28FyudTU
xDPEGbXCUnv7im9Rmsv2CSUMrbEe+JoomtLvfu6J56wcn7xJxgTtCu2Y4RAc345C
TPOMefcHuxSYYW/P+F4BTSwFyQ6sy02qPQlhBdKxIu7M6n7AE/YjuhEn3JGnwzSm
++7pa244nA/rnhWmMV4xMMhcnFs5i+RH6OKwCarvJd03GLTSCEOPigz/c9+hN1vo
CoNdCsU6zf8OgFM5DJwVXxY/DyrShyIw1+QkMVXgE1eboK1dFkhCikHl15nZPysD
L6HVzAIutBvdhm7Svx6IxucbTB81P4XhQHAbB0xZds02mogjX6jC2NC40NccYBy6
vHn04gG+9wviHsXarm5XCPXo9lXg4mb6wtwFWXqwWik6dcNihwrJ609RhLsAxWwb
Q/Z+eKuTvcbb6OYcor7bbg6Tdt0xLV6qfXssUjouxwwFoUDAz3ZA+VvsKuFW/yDh
DbLki7iALf42TIy9LFRbgA+JS2BPGsyIz/rfdcNLSlzcVNe9FmuN/58Avgp5osZ8
1GVpphQ660F0tkgv9Mw8+/zFWU9cUtaHnldW0cmgRWuxSAcuIwkNz6TclW60MQ/A
akWymuaIWYR9TDM74U+kVr/HGn2c4+wzWvrBXIKxTOloJdbaiv8HQcovS4jdtaiq
So1xGQEP7d6qxFFPF+0Hlpc/NwwfnbooSDTo/nkJAtse5THC4dHlE5dLiYdL6xKj
7Q8ff5SCoHGX8Z4jkc7I2rFLP1o1WAdg51+VkoMDlua35QdScccHHShqApiW4eco
mTAHubNQilOSSWKT4ZZEu696o/IqX2RiA/qwQuZ/XAuzsjRGnXyKE5IkzYNNrNEx
t/ifITme70BTk6AEd07RXNHw4ffpdISoP36xjjnWETK3hidW/s7fr+GqcrrqscCJ
oDvGGvu2zfb5/JpZ2PwQbj7XDMHsNj0/pzYu79M8c9k9HSTLyl/xt4xOGvsE6+e+
BO3YPPhJQGPS//GCYIXUyh2S/y68cmfGRqV8yNUhgDdhogbCgy4amNkZe2392RA7
xmyknwB3+pzN8BxZxJARj5cZIL9ijP9eXYMIrF9bVnCFYafbkdmU9o+iLQoX5nGO
cQ/lKbxXEbZmdYg6rr8EwoQzMwPLI5AVlE6zBETMSfCzbeoeXk/HZntLeCOZkCHq
uW1FSkhHFuGg87bFqKm7V5e0zSfjD9RSkF3AhqiEDEJPIG5qvy11p1RrH8CA9M1K
EfSk1R9ZMFDPnMPgcCDdDcFa7Vp9ZFaJtC0D2NKD9LL4lHvbfGp2xcP5rwklSXnM
lnhaTdQrjlV66Rp4+4OijFG9CX/TLf3jYvvuY69nA4/M1jeKIhHx268o5qZ0KaX+
NuL7AOjiHgJ9ZwISZarAleeRGHWheR14I6opJPq7/L1dtgJGzhGADmEZ6h43w+yw
kHo5jdTO77vOl2ZhtAW2RjSPJnhUthYSoKKmpAJcZuczzfQ1usK8Hf8EmxUEb+xi
fTQ5MYD/qtFsoECG4Qvi7WmKQNVqTdRs8epKtwbzxHhGyymUR58QKbbUZU0CWiVy
YbwZFWmuCzoDlAsfENlLUzDhxkR73rIsVMhH6rj79y5TqoLr2xJsO3yHdQdOijD/
nMHpTQUCX0lbhfbOSACCgDZ2Rdd0AoNBpYgiyUt7oOMHDRxSetOXjGe8jFsWVOLR
dN78ECz2QUSxQ635lbo3Np938W461hIuieraox9poluB7GeN59F4ZYyM0LNitRTc
Z2YNnU8luTXK1zZExB4Mh9x7FysZbhFVu3VJ1JudiUsZaZNobCoLXE0taHUEaBX9
WWh33p6JgGcq1/1sDoiHuSw03esCk18ILndoJc0lDMBXpNzKRVaFhkY9kvv5cYzq
QC5fr4BkZKBVLCP+cZrIV25x09Br44UmUQyxrELdIKILm/OtfrLucIpL1pEjUP5l
yv8uXoJXxPcJ4eUU9mClcb9osjkRIRuuTnEAEDjqnT97yTG94Je3WHjAeqJkpLLF
MJLME9l/8dpLYDLXHvF3xneOzJUu2YKM1Fe4rfVipF6BEbtIzaMCXQUZeGT/2COi
U6ztG49iKvfSHj0vf130hQoNmxqtabV9FqI485F7s9cfJYDnlCr4xiRfzzql1CVT
J24SSO0w/BFcJq7lU6i24C044rmNoIRGTR44wjpJwxfzMBAo5udPiOCVEQzFT/TI
i9ozinw7SIs7h2TRxWt/SNbUXOP6AeO6Iu6quFGhRIlSz/lcUWMSKpekQVi9hL6T
vfYQrbnHWhlToZR7YHkYawFO2xFK/ZvyWLUTRPfZVyRGyqnfmUBvxQRWkII/uynl
2hJ6jKjePPQTNPGLVZ6t1Lc+jbPMGrZ7REeJcknk90CvtHWfiJGd/rO54xAzJ3Hu
iaXFMUuHThRHmF1mLs4V946o82wunKvQuxJzOWXk5pKrkW+Kr3P8C19Xb3wX77FX
Gk5aoBeAZLsEnzq8WPp87GIudj8fTSgB0e1v1hPApJVZZicBizK/bgzp3Pm3IWkp
i8AjMgSNNjDX0tgk0sufmPhD+2t4gT8Xa9vTjCx1yzJo2GiAYb0QrtyZV4nsJPQo
ff6o7OeRJZmJBkJE+XDha+E5FrbCx/MrqKalGJ4bId5PUnsQB/7x5wsUifudqe5t
lDSRTWE4eJeARNirK4pXLSTYK0arM6QuCjAYF5yB0NGP1dsGot1sRZnk0Bpb8S2E
zddQBGXd/SdhJSdSNoeSpkoWcnQevVTDwRkFwudSTrDooRRAtdggErNSpAmp79Gh
YYgvDrkitxVyhPwcvS+ZWEwoZT6HZ3E5PzJ+auFpLvzZ+8D8G7brzZ4dEGj57XUF
76f+nQPGVu/ts5/lsqzyl1y4HmdiY+B0tgO1WRYpWKUb5kITHZitxoyEFh2QZHjw
+n5t6024kVv9vQ8YFBqxWzdEeKfFff4psyGfIJOFSGsrhuIOFm08W+HRJVvaySvc
pUx/e61Y6/7mb3Ku9QKatsJ2EhUcIqDb8CHH5yzXi4bfbd1L687JmV+2DDGmA6PI
SA/ZbuLVnp/8LH4Tr5Hqrr2NPKiMJML7SrPuccbjortG4Io4AvYxlY9BSthsqkEX
NBoiHn+3QQTxrRk5CfM+T5XkOOLORDXqmvSNghj11+MQZU1XujFb3LZ+B8IVq/1X
v6Avw4pLATBuVYpLOM0FdSVLsBuO9/mthLLq/OqsQHltlr1IQ0kc4hYuqGyKo9Kl
IMq1mnbX8BfjB95oh8ZQiWvr+fJOAM3Cz9W6Z9PNLgCpxZn32FyZVaKsQqtQad51
fZJkYqpDTH5JtMI1GaTtAFP+800rhQdLlBmG9VzZDrqCvCoLoVt+jqUGgZRn/sau
9WVqfU7aSfB3Vc7viZcaOLfKGAKLh9HpiwqaH25oQgMdoAXyikNZLDdC7wjL9zUC
u7wRzz6Y1xqYgZhSU5pSCvxadsjr2Kf9zMpzZGhtJ8GATz1Sr5dy9F+yZ4T+5evH
RzxlEj29EXf/LJqjtUgqLqFAD57IwPZrisHskcRXul+vriff2xRWAN9pCW8Jm7xo
bAne/oVtJia7v8V2nbyPEvBKingkOrLrTZJAwJTSU4D1Q6c7ZCtkmmEC6uBf8/mi
kXWZX492NbbKNQU89N0IvpVbCpaN+650xoviY6gVK3hUZC7s0BgGWS67NMnsTXhs
yLhtQtZHcRRD6W68YNR/jj4PtPSTCm3mU49/20ulvzqgmh9+zaCPjrSuQCwObWrN
D9RD7JkpI7vvblQHFMFMPYe+syRF6XY+vkkO07VR++pvsy0LPsGsHsz1KL1xYoVu
KtEGrqOY5AM9/As0Hsv5nXVQQdEpUrRyMIT607jy2JaBGgxRNK7ruic6JM8v1zga
tIBL8dTHY59JHgsvVbxpQ/uExwXbkMFn84WR+mStREkIqztrqMvE8nY1Rytxw6OK
GFtqShukvWR+fLkhEL2yIVO4WOnVrynp0i8lNhnMnINu9paCQO9IDbAON0AG48cT
HK7v02vTMAa5y+soZ+1TOWJh4l2s1OKYgGB6jqJ1XSE+xqwQjuIjBiOwSJSdDZQb
3sOSBbe039CCZVmIDMu6d8gKTL2zPLGdwmR635oGdPjlbMaOfDAP7ZQgW35AfSgD
A/IKZaaxsYUZ0mLK4SGkwJkZPhbtBM/Q39Z0jZZWXcF8conRcPaPoW/ua0Pmb1Pr
1rO87j8FvMri4mSrxhUAnvoMcl5A9k5oJehK9m/Dm+umvsONrvJvf4t05qmWdnII
XBdtUlHFXMJdRAvL0a9V0x1mLww9Bcsfd6GLckDJOyT16Qm562yjbr75gy3itfAT
fDaLR7X+3l0j2pkdOcN79ZonQGY5+FcNJ8SvkNOoyaTbiTDNB6f/YDwtWfe1rZ/S
vnBmox5TYL52tj6J9KMQVk4avIYwq3X8xD0jNvfX8mi2idVVVAR8KL1EZxB6g0dx
z7dPNEn3GvCjIYJK2Eo/KLynyWXx0U9p1g4NADIjGkIdBCfHAtJGYvRZRcKsjVZX
0DmahwSeV5t/estj2I5fL1LeIzffLTmpLZwFSrRNhsaAwlUJCti/H8xBR2QIgVjp
sf2+vrFkTMYigRZWmsJYB3AeYevzN+p/Fr6ZxB4otxXInqk5BBT3ZSuTaiwzTOSP
N9OdjEKqyi4sdunPElgvQo7rsmINx3Kt/VcEbAx/8E1RoTAsp+rD/0krumMxipV8
pXmcoGg8aA6w4MrI9LM0vlXu/fKZ9xJtWH/kmCn4+PNljoBHHqGs46ganVTPN8Da
eLNenPv3WzXYIRgtxHTh7ogUIBP6z4UCRQe24oxTULwFgCSY4K5TbC/Bqyp3R7ns
+/pHFnECYiAwiy3385N8sMKObIZH5ivW4MV00fYamTrlywjUxjQz0ztUHvkT4CjC
lfXp039WM9bk1OWI9bTxeqx5bFQet3thS0gMRLjLTmmGt6HAsBw93b6IWMqXr3cB
kOXhlmqtNklN2ZYHkknI6l8C8QkYB656PU2miT9HbqfAFKkp5qBaUxyuEn5L68Qv
NhH8NTIYv9eGArn0BQHHvJbWIYlbWPup/364DLQPgr5xUqdUpK0VPAJo21hqB6cw
GTIFZ23Lr9D3Cqu+aXw7iSoN29fdKI3zrbcAcqaUrHKAQ/2aEA1PBYB6qqnNxJTJ
eKj1fubOyOJHU0J1Jw/mVd++imHuEyoj43LI86gkh/SDGAoWEp4Il/NGN5MeXEyB
TOmfbguloI4sY6xtPY1EXdk3sGmTDrv1sI4581TU5VgnXD1ieI/Vn2X40OSSLf9I
t71fWfSP6c6Jj6OaC84gSdq2yYrpIgUbcJx1UCK5ygH94u8JLgvJM4rG2efHjhoM
uo9HQNjWVbFD9ikKbL1ZJPN4GHUXyEH/27Eg2ZNSyn6FPIpivWiiiQIBqhU7KnZW
fS2MTBmD2I1OYxy6KTTcFpJJxuz3VQa5yiIGbgw66RxBXqEaawU3BGJS880LUYi2
0ZiKn53qvX+7YHYJ8pLKjISUIbMz++x1TBlmkexWDGeUduVcyhMdlYf/C+2w51Cc
8RtSO+ATzjuSC5J+JB/Cf6GqyA0tQUFqPCVA01QvTBrlWANdG0547h/205zIZM3D
Nf4yuujWjXIoA5pL58Q55RvN9ezvxK/G+A5Zm34jyy2ks6A8/afANh9NCxkiBTdD
N324Axil97nlCVziYitHPUeWmWLS3DEXuixBnqQp28ug1v1EB5Dd9ffWnMgN8yN7
0XYei2c8pwwxnutTc/Ef97JkeSsxK/+/5ENlnpHll5yN1gp26xsVQQlBb4nSffnz
gIbTWyjA0OaPYRfPIgvuN2sNE5xKsrkknF3oYj70UaL0cXkMmBobhiHV3soDNI6+
7G8xpO9uVypnOivw3L537soP9eNLBj2cuDvJauhRAmmU23BGb3e1nu2T/09M7QOQ
m7ZXuMMdCoBLXW5cYaGNvOPGETU5P8ASVRh0WPDIXk9Wcppl+6/95199oGLjrDXm
8+S2zEC8fJRd5gsdpdVyCIybTybNwar4wE51RsmS7rR/lTXDlel+mdjPLgeI1Jyy
/hs3aGT4Ya9jAMJAAbdiV+291KQW5Jitdb89J0bnnoOn9Ozx2MvDo/D2YHfRuDUO
Z45q77mfoqOL6USbkI4IqcpkNFgYNK3eRL2Gfuqd96QR8Pe4rrk/M6gbHzhaqkbA
Xe6X4vMl5WuO4r6iHkpEQBWYbU1///eZlqou3TDOPy5KNINeZnFB5roda5/prIQF
acDHklZfWVSo9/badGPe/jlRLY26SbMfW2hGX1oJLsHPI2l31cqFjBrbDzaNCpY6
L5Rq8Q2ggrW8Ca2Y2hKxt59Vu8GgVhvsvya4mfBpzw9fUe7TmO0TefHtm8m2qxtE
WnBaMhXtZeHCvHOSQIS6fJoLmJ6yIYU6wgtp4v8P8zctSLHOzOyg8vayHsHFh1Zk
iT1go7wSImniZ56XD+NCqdZz8CNYlcBFChug+nrVtvUTPWqmBqLLbxi7TxWkXGI5
HVakikW6dRUdf4brz7jK812m1QhcJFtLpzbG8ham9c6c//uoCCq/+nm7xKaHZ7wh
jDwn/gwvOfvjElqD6RWkqT7BtX4Rk3cAuy3tTMtFh+hc6hOqIMnzQY1n5RBlXq7u
DDaRHc+0mnODDtE87oqeRn0bttPMq2FPlPOpzj219KL7yVLSLmSE1vUN1MH6ZCti
eeIyIHGV6kZ5i0UIYuMQ083y7JB0JYlAXwpcnQx3dY3OepSUHPLfFcdNt7/9shA9
PIaCk6382yK4kqKQQZ4Kf3zi91SV/14ug6lAMw8W+DNWQV9ybmpNu/9TXZIxqkL6
SIZGXMHkpH+BUcS/gk1FoJDeZ2pL2r3JuvrAlFqIjNyc4LzKlXe576zI/P5tKFCh
A9AA3dK9MhU4MyO4O7YPX7cclL8x7lsAhChjCHBYVkOH3/UjzUu5LZgXvA7obet9
AJzYnERlfUcIHuFQfY1+lCbYojCdQ1NwDSI+7ZNLpm14G45LIwGBH5wuwSlUXc54
9ovpadZB+hTgOlOKXdlvwzkADTPeWAclSFXRwMQTqpEEEY+O3AdBV0Ye+ciy3FNj
KUxEwmjrSMbi0eNDaHF3RqZozOZ9pX43yrW9RvbZZ+YaZua9YB8ndwurDJf9ng/B
BZe7mIBtV4pBELRnT7Mpz12RDC/lYUnMiuiiRe7Q3rw5g0+rXuxvKac6IA35ok7Y
qEiFwzx1zGEjyvQw60U9pS5MZAh/t7+Yau4TXutgsIAEBkqHPA1BurPfXF8R4X+3
psGD46HWAwwoEyyZLKwQ+kPt7ZsLx+vPf0rSjDCiEvXYxOPLa7jrVBIvyV+GQZcu
kkcSJKNPf8Djl7hPRgTiPf4WLS9ePl+5SlZQ5bnsFqN7+9dawkywdDHPiNCY5ghq
VG0hKPKcJX+8Yt/q/PPMFzqOn5xuB5PBG5qL4NDCW2OyRhdnB9Qh21X+C5U8F96E
oqyAVhGdXIgwX3TgCYzKH9gQNEUpfrHBRnn9v6Q7nKeynh3X6dF/Pax4WENZnxuE
AWUSsAFdqLWWreSt0Af2kkeWwVgaiJaYoEbLnBNGeeMWW712Kk5JU67pbyI26I9c
aPFzFMinV5f+o1ClAFH8V7mfDi4E2z3SEiPWPY6cYuI9Uk7Kuy9f3vRy9r0n5zdg
D0MwrOh1OhJ2iO4NpyoJ3iNkuKGrhVaUhVP1vtH29/85VKlFMcJ9U1USaHlzodxC
oKVJQcxA0R3vcKneHXYldngLrN5/pIGEJPOavu4X3qGDIwPdrHs2WjkP+u5t5SLw
khHr4s1zs9tE1aJhIWP5cNAtwtYF3n/jAG0THOMHRrr383UibRRzsyBQDHtoTc3T
aRpu8WN0S57Y6qgATiIOZnd2+8mLwD75DXaPna0BOC6fbmk/bPuggUHNr1Q8u9qK
Og0NAuQERxKhfnj0TuQPqpVIh/HswqfdZQILBJ7NJ0G8uvPVFiVTzw/tq8p89hbC
cfQ+j4wwAjx3cL3kMHXBMRUphFFHO626xRqCcxdiWBSHKrbLejEXJZK8SX8uTXPw
dRW71QRFll0rUZtm6/ttSda/ZVluVG4G5ZWrLbQpF+0pkDYFdax34ITZoeoqx4jd
Q8GwcAacE4zLBaPuvPREl0SqTkPq4F/r1PSZKPIR3hhM9hWh9Bg6Bq9fvyNQpH7j
P5DzMHhZHLvtn/oUf2hLSDc4gjR4PnqH2flkmOK1BH9Tqe90X8eEmJExA1vi12pM
YdOzcGXL1bQqbGJg5T3GVJTgIL0xPoGw5a72QnmVqsAiprKqjYBnjbujxbGyQAuw
da1Ek+tMFGRymtF40LzL4vVObLAY7mJFGT8q0gbYaqDj8eyD1Mgwj71DcxG/fCSk
OTVJ6xnz4waSMvf/jbMV/dhqzyHT0T5VVcCd7ugrgazCgTaLF+YWe/ICdmFGb62p
NDIO9pNC248VlhDxDmvapiHoprt+wfUj8o0EjJf1uxclgUmmNfAUbRVaqdPuerwZ
dihP26x8IsdcFqCSq76I2y9gogMp0fKMex082+2ojxkA1pBtYeNODzzpIKAgYN3F
kfQChFBqIpQmcK02JYXfkONQH01d8ieccYv9q5Y0X1YaMq7gx9EUedqNekHk7shh
lZhrTwXsOS2UDYtACWCMTogG1cuGMvmftQuGDlZ9AsNw6omjIWbAu463qbNkJ2lT
T14x868xS8iljva43C/8tJm07ZeOIIzIpml9RtvvXfNNxAsGXBeuHAy+jwrC1GVS
2qVRj5678n+bc3vvwQVYauHJFk+6r6MEBUViz56XbPFWrzj6QNRti5suK2LsX8B9
pEAFRhaYNF+2u8N28WsowgtirVDz5Wr+UyreRGuP9wvLos7Qjo5VD72YzZtCuBDx
jYatbBRoD1SpV8Ar81QMKS5yhp15wjrqQq08qGY5uRVKqHg4BynAIpdy0AUMhllB
1rrqtyh4CW1tH2b8EdFaofZkOjuhH6Dc1q470rZcL77A9aRHJU/NJ2cjQndJMEjY
dmq4NvwSSFtYfcqHuDc9anWDVrpU7DmWq/w/iwDLjTrjmejmUEnCzvaQQuNVINz0
WI9Is8zbv4X6in1jjpsRWlvxn+/gooOYEunXLDHSmI/9bbEQlTS9aH85L2gU4jTy
lvNF6ZEdohlj6SIU8RXYUpELy1zYvdCICxzVeS91ATGT+nq3o6HCot3fFMj8A4LI
RNZ6I57x9lCVregzUcvyvo1aypilJWFMwdN6dYYMmoJ+85P9rkA+XFmLo796Lmgl
RX+UhC5jin0BQEFUdNCJddpOEykg+q/F3Rt6KQjdqN4HETNHFX0foglVigR4IkO4
AoIDI0YQc9jCal3cavcn85oYFAZ280L/k5WR7SruK05aeKXYAZjfcoX4bwtk/rFh
RrXy9zpuTbUrwO4XqIaIm65czvDhUNeh375kSC0S2sLfTIGTwWxvwdFr8L+dAHxD
b1CVNnqsRLGNc+n+78cz6BWZlpMfK5zzLWKYKqjPqmOof5NnD04odq+kcx7m6gfR
aINf+ZaCNSdaFOC2mgcoqgIxvDHyDLL08Ce/1s/+KbGsUUZJ+Mp4ToQeLnBgXyX8
d8wfOxDMngsvaW0SugR+tKMBKMUuzLNT5/3/T9blNFNCIyoCdYTjqfugwx3n+jer
U2I3d4aVLnydeJbf+Jp5Ks/Ye/iCG2Bu6q0nAWc+EF1Oy+ebvWcoJ0XbWSM/MnOX
VtNFauJsRR4Izyob+XL4R1F37nKONNp2AKZMjVoxnj6kVp4+YmK4NcLyz1UOd8g8
nh482+GGmauPD8IOLDU3cWpEhczo/JqNwWE5djppCKkbp7asK49sQZm6aixBVqbM
Wzp6/cucyxiNatnvSc8gaWVhGFxB4SVEIyqyncbzS6EK63F9qgs/Y7yMgYDVfras
2bKkqchlXyY3fy+s9/QSHHdEGjV1PmOWAt5NGSSrGFnlb0NNRK3O07FBtDBtNffx
y4SRhldSCXhdMlTOP5hKdqBgBDp7RTsKXxEVJUYNsJCjU8NeXxh5OKj5dtReBrnD
y9EM13zcOxX+DwaPJX+va+hiiGi8iVjszerpXhVcdeL/CCHqRJYhxzio0VroOA+A
25pS8945DlddtuuhSU81mixE45dftWZlrXTZU+40M8Q2Yi4p155d/zii4kznPTUM
htkDD+Raz6jEeWnxYm0Xtpj+yDbtg6zqP+ssbJd6BK9Y65tVEfJO13kubuQd0cmN
Ifja9IMlk/XuY0OjLHQp6tEKq0KDYEGZiShn+TV9S+2IxDNdtVvct/vFghz2WmeK
iJfYnBr78ja9yIn9UKgYV3CtY0djwMEY1ibNRIKYpY7VeNTau+5YBP8JJaYaM+2C
OPT0s7DsHzQrlGw8CGMEonnr8eGZqOSHHVyxyCdatnn6xevr2ZrIk3WICwjWneBy
MGICn0vtDNjjJmnqbKXTku3mjqZuST6Iap7hWnDTyyUrZWsbBxNKN5ckxb/wciSh
HPMDOGkGyCLZDNUQPGzDiQF9Q7ZoXHRoYg9/OL+vlxYjpquaCK0qbDVfTpNMYL1w
5joCQDh0RGf7YEPRKijvnq6sPQ6QqH8kyzqcAWynrWeGe9UcSmB7tYiQcwQuafnt
tVAdz5TvalgyM2OU3dC3Wiup5uqCDMgEShgoSIHuWWUYZWdJKBGVEtCjDZNhmIvk
UcRRbgRPEn48+ijrjq+giUs48vB1vZeTNO0yeOK0HzMWw/SQZUPPYUtRSk2CSSkC
syqrpzD6znT6XF1uB51tJDwxrkRIbziROP9U0MbAxT0dq4nPKSEDJS3WldhLhGBg
aNbBC/hbJx4qEA8FYtuXZj03d0Yq9X0HND2t0r0gh/LJFf2v582py3RMmF+f1NRS
l3AdVXiRdWP8vvs/TJTewB6qn4Wp8jQ10yg/8pdYC0xgBkaghypNWJw7XsDlf4ui
PkhyKK7WBoXpXLhmqNWXvxGawDPxY5UZbnYowQUztldmow2NbaJCG5YiGsZVPFld
NEY38txrzxqYvanLJbWrxq/TcF/NjmDNAMInsrzyTJltQarzXsosVGoNH2WWAF8O
TT1k9WqRLAF5K53Em1KStF3HboZGHx3QVOmhFIAulUmTce1gQREU1ZyRmuw4XnnN
JFmbZehFNmx2rf+67MQHXe6JQmV0JuZ4dIwyxblz5R5xxanQwrBXsb5/GEPCKWrW
fHl7pHeOQpJOfNGpGibGNTWKJp2hhRvOjnaqmOLI84DUAF5BW909g26rrF3aGAh/
hynREXQ9DQ3pMFx83ojIsZfuch+fpDc4K+Tr4xoX9+u/OMQDxUZaY8+o7vugzAYm
UHlLVy4ZiBikNNeY/pppxoTKs+jpLGrauFaMdtTgMxKVXhkkiXsMl4Rh5j6H7tAI
S0iFLTLemEilQSqAiFuLpQbXdkp7Ge5Os9Lh8byPNO0GIAL71rdW3D8V7fZQKk5D
VGWimVgR7RwdoUaMxC7yONtPTtUZhE9PTe3AjFhpTwOCEwrID9WvI+18AHA4Ok/9
2CrWrmxNG/EyGupKso0O1VWSG5zpbxpY0XLWpUVaD0tqIF66ogioJOSj4fkEaX9d
btuak2c2EnqfYq/f0fpLUSIIZ8ypQ3KWvalk+VkEFzh5d2Q9vKfLCS+ll9s7cmwD
DDAbJe5zwBjBB758FkB5G0moolv+xBZNv7mwKLtDWijD+CHV10tuHISK2wJ4gM+d
Te+nO3YdjOdQMNZAsz0Sz9etZYCYaciBCTSJjxsc6RtUkGpge1j1JjoVVkGHBJpu
0tTyAFMxEBOyzuthQm8KIZlSGmHJ0FjNXLY9bnHPsj9mqZpKE4UF8x/H24Zg/W1/
vKgu8bDbOSh7OEqgsUZxMN5a0EnQjs++hmYDtmyJb95CC39H1r19ztRGl9lsphFp
ECkYwXVTaecoKlBG6KuKcpdyH1n8WRTdKG4niG4Rn2jpsXIASblOqJSOTHJL+hCM
2beWVlY1ErupwnHqmJ9hvuyqf0Mwwgs49mPCfgBA9DQk6hDDjln4mXqNb7+5mEP1
+23+VTxKGyd9aGjV8eC6NsfIXPK91HKlTNxeO3Tc8IISfNpeJQGX1Be36NzX9XCx
ryN+F7hIdR1937/CbjT4lT2odR38SFUMkeg0gd7nzXumhOFf+wfLidYCCQgDqe3j
LvHM0MlLkc2zQ3PNW3Fx36IQlMpBU5QHbjM1RFGeF5pmbAXkmFLly2iJX4LrE6NZ
SefOMFX1fHDf/MLaDpzMapfzFYj9epG+XN8hBdQ4kGvgmApW/usewimXvlN3qWFk
RrhKFJWAm8gBf3wNdfLtnv2w3OeL6KLZbPJiAL6DuQRn5itXwsF4SMX9JPegla6H
M1vti9SfhHD5eKEVhqLn2uhQe/pDTUYyWXRXh8v9iFpgq0Mes5xDLyjV8hgnNjss
4A8AnrEf1SoWpmiq6g1XyUknrmLNgvIfFM4v3Qylm6V2uNqJOLxoLOgXwP6JI02D
z3WOKsr0XMLyFQ7dTQ2Xv4LUwkISjsbJFTxQYKadavjyTsT6JDg8h01/RfurokRY
y7Vf1KVkl/6hBpGbcWIgddSDTS66p94ULXhnZlvb8y9h+eyDI8dCETj6vBQ8d+k1
we091zOBVy/ZnovtaOPUXzBYNJMQFBoRAkQpKk43eTFjwOsrsZkdrZm4mV0nhkqb
a9MPUNl0/pSXJ+c/toq3J73nexmkhtGMBwrsexSElXgkpQU9Z50BYZY9M2A4ICtu
EWC/r3195fcERTFiN0/yqvEEojwYvTEaAGVxIPfP8UcREfO0SkEyVQNEhrITxEZK
RHIOilXpeWYJW6O0g5flGTMgKVPfqkiWlz5l+E4qoXZZw0dJlPmo4fDmeSIa9st0
HWjIRvF22CDS3Yh/MqCotzHDtyYWgY8auk1jmmn25byDLVO9BVUhcR11ARdK4FwO
gzhFV4hDexOVzQM0naOALtdNf2OHbeCyzP2w5rgVzQOahaO/fk1xQi/Q8hjEBOmy
BoFy77KGCI6Cy967zJFkQmelGOs+0/Fc44f9lVvqdv01GEaw3rN6WX+iWTxUNEow
6Xofj4XPAm3i4nbsSJ9nb2c3Vu+RFwr4QsxVizyrA/AXMsVu2CqZ/CBvdFdma7Xg
aqBRdB++k9JjFKKs5C1/0ajyZE0RTZ6Ef5CNbS3B0T6CgrDZHxFxLdcADax58Xte
wUnImTFE6GYQ5BI5kfxgqiof8byfmyssDrMfPwjcFXGi0jBF5n4AUWpEI99Yi8zu
X74VZ0mvtp3MOm4HURAfpKB3mTK510BHUWIZAqLmZWJe7NpAYFKYntxoqxAXjPap
x9yHhKAQNTAok3hOwiK5ps0rxYHGMoVopBouCOMt67a2G3vBe8lw54433xswyMpX
lL4u8xYZCj8rzyUZssYGj6mnOwHerW/TUx5GTg4LeP8Q1VpWxB4vxPLFcjHI/G+7
gNhauM/fqBiK6nhAYj054U0OLBDmr8C9o/kHjP9oeO2yIeVsN52h38rEuP36F6+Y
Yf0WpS4sLJf8Z3hQbMaWng5wEIRLkIOM6Mcx5wqAqlwQJ9Sl24p28/6qbQT/IChY
HVzPRQ6DIvzi+2wZ/19NllSl40uDcLjufpoXO9PN2YPVjS+vehX6PfsZY1u/EaRX
1aWPLmcCI3pDdjTtM6W2L4D+ioRTUjQ0wLlW3NdSHJEFjLqXnsL4OTqUSI+H1K2F
UZgR3N0HCvPIZOciP78UYzYzDjW6OOFxoZN9mj2fdfIJS5TB/SLRTn334X5UfXQC
FLg+f/2cTpzSTW3P9t3GXGrKvBwx9o6nTGHu0vjTW1HDFFlCZ6YU0cEbNS+XbQXY
5ZsOmZHLZFzQC6I7JSolsKt3J3kOu4JQUaToPr4j7bJ9UJTaYz1zNodgxiESIYpg
7PyhfJYJLk7GK8SDFhewDD0+sbYY9bELfCv2UlmEtsM7pNix7jbJO6v6rn4lO9HJ
I5szq+cXY09qEntyRIynUZ3czo3SQ7pK6GQ6QUlIapepaewwzQYJG9ihneHm9XJ/
TybvbI9zJjvATC3LAlPxP3xW1lOstUU3yjqCMqugPRFdRDhuF35DKyDnrP9omaZ1
cp9bSDtdI3YUoIwP+/qgcgnz7LSxdYa+pSmi6beY+O4vIIFuizT0H5RTFX9ccNSe
uco75p1QNa4xmiPjbqqY/ikeovYBvVB6F2OwLKmTRyDNjlVcS2/DzyH+gzb27AkD
usapnL5zqnz1CcS44LqLlagFW+KCU0RTuVWdkyEz6wPchmJut4ZUsbyoKnrlLvZx
tMkD+180bdM4ep2L2UCVMou05djJ69oT2D+/Q7xnCXDg3sw03A48SFhsXemvzcT/
xw+q9e8VfUt9YKQaPpgNASpy6V1ftHcWFDmylX3u91iAPHo++xz2VSrVKsMooRrL
JZniaWhQhaUWo+Nd4Z+eKpRmvDmi0F0aLxzfXqokxRsyyN0nP9Qcj2QJDwij9YEW
RSSvmyNhbVO629QbvI8JODOPK6EXmEoxI1Hp7tawSE2/3wuaZtkVpAsboC4colog
MNs4yeaHZU7ygSm789wDkX1OXlcVlOhCNCvG+mXpdClY99bgEJQdJAjQCRTavULG
iCzw7n90RoE+0IyHfSyup1TotH2vQd8Xv7NPmMoc7aaf9IUw8ooDL63CTFr/gcyW
6a1gb9HW3xUrWFA+mM60QpF3KBXTrkDutPJnLXpD62dR5Fr/uEuGVHuJWANGQw6x
hNo4V+oBtI2gmCwMTYMi52MW8/wrHABYUB5uiTcbXxsuTVcb6bNRKCEQp74XBc/d
HW0ZgPWsNXVE+2dACW6/mDHjLWdw7s87sIkV2Q9VWZGAwBESiFXFYiQ4b+znD4VJ
U9LcLvu05oaG2dRBOvqFmkFnJF5hXQvAOfZtCXdfgfw5NbP8QxDG4oHEkNvXzg6o
nKB1D1JqOs8TqvB9B5wz302vzHaHZbFma71j8vy/Y8ZOlGBgYUEjTlwO3s4nS2b5
ONnVqxjuMgAwraw6reNKXEyUGw5IWOUGI0krWrpOGiB3+Z9c7EhmJDJGUy57eGHs
jpxRRBdHN8WR+RlQjlNvuLDN+0CPbLUZWhLBYx3Nj/IZeHM6+zGqAUVr5lfZuKmM
Fe7Dy6vPMa1TPbJqffVOB9gffVDGmwQL7JcgW/k+ZrjN0bCPajnRte93Ga+Jn/RV
VA5RGxtFkUBNSv5dhgaipNsyz90Lv2gIhOzMD44lBY0rLt1ttj1u+q3PuiDc9v6K
OHO7SA0xyXy6I1dmEs71nRtBP6mV7fp+M3S2CeLsx+78YJcfpOmKNO7ASI7HpsrJ
komWOajid1tgTixA4f9aSDJPAWwl50nuexb8X8dcADSLfv5sYfHg2b20slhTaOnv
eVYG4V9rU7oGyUiyMyR2hvCQl1lcqkIfFuHGbjDsrNlyMc1ZeuoFL7y9VWa3fd2f
PnD6NgxR/cU5R3cpA3DPniDhZ7kDP4yI4aIGxR66htGZsaiPODj6NTtDgVsJZ2Jz
ifQpGBtz4OmjggAJs/57+GRrGtUwjWAxn3x6r05AjGOKaw2OIpqCqpR5rGskEq7+
QCZCQjgMcct3EJEsHp8e9H5yjFVe75jI20qv7qF3M24s4H+p1q6AO9q0nzrTvFLC
tcHCU1pWLQGEkWOVeCYfqsfqk7rPqyOcUfHNaD349IGfH2jxrcHHtxGBB9kmCZLi
YN2yaZJU/V3fi16gIRDO8psoDENdzY6eMK/nJb9utqMejE9FgL8LpzjkNYKJ5blo
vjmZHlQ04HwSHaZ7AO+GCsnhD63ahllQbobfz5AdWQn3+ueZ2WkIacJWZhlBCVxe
tS9TH6Io24ErvsXyGF9UGNgtVBAKHlbNqc8SQSphIUO+7Oc6YR2fkdBJpL3ZiwJO
BsHA9nSPNjzLiug9WuLDB02ryAr50WlLX253FeNSZax87DHEQ+i2JCuoVKntkc+i
SrBJziPLsRc7IxUAoShH6765QavZLrra3U1OyAycDkqmeb6n2vh4oWApjs2tN0cm
RuXS8kn4Nhl5A32R9aCW/+C+rtUxdp4n+VZs/D6G1L9OP71wzqGUJWvhPnMj88og
WInV+XNvMKpj+RZNd1+olpNQQwAmZPMD9pyFtgzJPfm+5CCR8rxOgnY7HCQe8Egf
xN2gsdAz6QAQmdEymRolR/BWE0XOuEigmU1gz0QR5g5DJMm36z9aAk6vRtKMBjjL
YTPbSWiX6KN0Rs0tIOl/Dkt7Yu8tv0IO6bXdmpgfweMGmXI9IzRh7ifiAz7O2MMT
g1VSgUwOi3T8MbMpsgfXE/5SPRpsGyaxSZvc29Y2IRyy92cSn+UHzheijPKkzzUx
K0oZbBlye09ez6P8RrC3zM/wAhgXFwOopmmJq74MjDFJcCqse+bT2gTjXAGwC8gv
z/D3CW5qVI9rMH1VIFaifmh0LVwIhqV550BUu9M+zz3OdF+e5wNdJ5nRulJvV+70
JAWyYXvLfwKeCFMQEL5DRugiM+BkRqX044fH8JgtgLPabkFp3pXtNxM/5qFUkxwC
w4qWUaBfhME+1HZ9DXq3aCDdGkSMiVW4TYpG2b4+0VMZoV/184ObFuegxW6e3wNy
zhb4W2P0OoqwkDEoFrxyiiXM1iqCNVWKEtelQzZL6nmyKpBcpsUYQzLxwJ1jv+UM
oneuh2lKMF9RaaIXxe8O5Hb5Ry/vjkpiItuvBllxalObvyvJDgRBSmqX+GiULREn
ORjcEwYUSM2Cphk5TzWdA5zVoXhNVY+MKmsR/r61Uxdyv/iot0QTOOr6GTaMu3xl
rUABmXZtbPX/SxctegVkyR7By9eviBLUMEM361mMZVsMJWDn7mpBMnEZX3YIaDl4
KFar61JQa9tqVQZB+ee/nuW5GHT9Wd6bA0v3w7PkDGdKkaPjSorIDqBFzXR95p8y
8jD5PaOGzu5mUYJaXqy/BU83N6Bvj0XulaE0lkHj31N+F3bsP865LnzuGVJ35elU
3vkvt5Pt9vQ76khRuZrT2U3pnvz+7MyORZKdI7cG5gEOPczuEREVgbMtkGhCo+hj
k+lbrMeUkKyyjUpd+scKGcP6ZsSlgJIijWB/P3XxQzaOXQ1bGmR0MefwKWGKbYtH
x9Y80+7IblyXT+Orj/D8L5QQXCHg2hF7T9ujGtjwR4oHGltD9rVm1kgMysZt3TgD
lHUJnCUlWwgrnXjwXq/iRSPqqCzAWcVU3mmUXwDAz7iwkwag4Csp3FCjCHZhzjxF
ffvY2r7gqBX62o/HaBPdQ9DiGjSeYCE5neMo3p9mOCJp1bozBFp0/p3e3qRYdLM8
0J4su2GQ9Z1B5wK26mw1qL8iQvcuvjf4sKqvLlhovjpslJcQYJjAmTSc8iE/MDLM
Fg2rygHo9oH9QFfcVSPLEtRzEyQRCIYV1DTPvj1AF+Is16N0cCqIYFizO+HVLJ1H
vpBJNkx66Pjo3fFOrJXWhX4T2vu7p4zBzWf3N8ju7o7X4KQc2l/d4tcmonVqszog
kevHMKQXGb8i39woQ5m2TeHn1LPIKpotAMh7rrHmmNNrdPuScygaSIE9jsVk1Mrk
2v/QvN/N0W3TPqZzX4uIgv0e030InqGkV3BcXPYqog83cad9+kwGMrrn4XnpRrrx
82Te9t3Z/4OnKjRDl6FmOCjm88PfwWV4ndcm8KqoifmuZO8yUzppZNJtcY/SKjV4
bhk80Z4W0EO+GgsBtfEmBQb/h+8lOzohNHvsiU20mPnfMXK7B+v424OFjYfORhVl
pzMXciNIPcm0MecnJ8G9bbd7dohduVy71fOH07FlLifAM8mQcb8lePIEUhdKdrAp
54x2F9VOUzvdV1buVvyvrzxL6zXMxXhFNMKaCgQd336mf/X1wusEOGmqqN+I1c3N
IChPghnSkuaTy8b2gCBMnD19cHvRkQgBpQsjTKawUIpzeD4Mvb2ZGxtWfHOKFbH5
Rz9YS45C9dUX1BGep8kgyGleZ/q8Ewc32ogwEhyhWWBfC0kUF/UfU3F81ek3LmxR
dyJHcYNhUOcYGhBPTIBoTpKeZOmDS3ZkPxlFUXzmT8FIzK0BC3BwHBKE2Qf0V61m
VFYH5iTv7siPW3ZPMrEPg0tztPjeActAJUmWlMTpBfuch0QxN5hFs6E5Tcj4jt53
x2BajA0eKWPjVBY7NEN8su1aP9X6ifmbcKrS5+wwUygmgvKInQKiIgqz48LoQIrZ
h3tFrwmY8qpA6F6IkUwF52O0EDFKl4yGgi5GOUdmkZffxgxfrB3OyzA2iVUu0cng
lWZ4POxbQsXWxNrr/Vev6j9ADPn0n6Zbq5hp6Q2grQrnGnX3qjYs5E7czZ8Apv6t
PAbQ6w7tXWuUPMjypm5ZfN4WxcwewPWzefpEl0w6fUHvmPJl/EClAaj/GsomRgHI
wM990emdLsCkClDqvNF1KxnD+SdOhPzePQtGS/0F2Jxjwjp5ThS8eFix63aBAuH2
pGGXctrqjl1pQiCLU4J5IKj/c0N7zsxqL7Ts3nlYsluhEy/NRKl3pLvbQX/6xARf
c8grqpbQoKmt21NL3DhKfvJWZFTuQNKMvcVNjTkcX8UIGRWL7kuOcNNLhkUJSPuZ
3qvRGwnqN7f6fGDFLJfPkH0sSVw4VypWN0GlVeiwC1EyQJW1t3CZ9b6JXtSI8sW7
el8AmyG9dCLEF2efQTSMsDjHV3ENJKlPafl9kReL1lrSBKxxinQWjMWb2Kyaaw0D
mzKKlJ1e8n+UASBui8OkmvoyBiv4p7CyTJ29rjiDwYjcsvt3iBrxIwBSXhfJgQN+
UaRVf2AlcuDeZXoKALXfmGhpk7M4rVskUWjMHRJdpQM3wXd57yx3FMsxDExTO3Eu
tv1PEQmnIu/xtvxzhFwZOMFDlXctvSKak4zKHJVNrVjAcVTp06eXc28Ip6GuI/bQ
jHrXdawQGf5KBdk1wqBjE3NhQo36qlhtgGFX12Ifja2tpm0moLX1yI3wZZMMrvTi
v0LMEEmfUXqlkMRJ4LXOqxiWqzK19XRZMKUQaEOqY+HsW99F1692Q+cYYjLI3U5u
I3i6LoT6wOb8A4NH/2yuyxk4QGcptWqXh5IsKDBXtlapTssMVHun2tXfW/CHeo4V
yLEf9WoyauYxQPLRDmdaE9Bayxd0xmBxpM6wsF8jF1ZD9ZweWFRY7eo6iOnvhOJo
cHpKe4A3T4H/TKX75J6J2eeRBWQonGOQ54xvneF8KVDTFYS1MGu+hSSkFCfAf2ZO
UJJYUS+dR3ph1RkzMuPzCGODPfrZXdaRXaYdnorR0pE=
`protect END_PROTECTED
