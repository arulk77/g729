`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
gJUyAxnJi7CR4KB2qfxBastEc5tW0/QUQ7kKP8cUvoeT8BehFKNOVPkqNL5TsNAH
u24KVHnHkuwDUinP3MvHdih955IMZwNOrcuO/9376j3MPrYzXEKzzE3MjO7nyR/k
C4QX3m0H0Na1yeulUGny2szkMXAHMCS6Db3F5IVKW6DYG9nZhIVAghlDU056yxYO
P3wZBh05TT6cXwGpevL0q4y6qOEgot7EBR0vxOgrjmSpqxCynu9dHCUI2vn/j5mn
dbFwwY/vkzUxCfhefYpNL7yPAeRu/bF53EYJtGS3FYYYi1E90HwV1bsCrHpXy1pV
H4IYBs5/iD17FH6HEijclggQ0KuJxmXYItm3qkRsiVs=
`protect END_PROTECTED
