`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL4FI0CKiCodVXtjGAvywBZLggJ2jRJTGdfaw0XviB4s
wNyfbky3kAX1HbwtNeW6CwzopWEh5L9ieI3U0qcCynBqlUgQdI7xjqZI7v/srEbk
XuZH21UPjZL9d0Q38XdINztJfj6SFnY08ymiR13skzqUpdFvaUKHtmHCBgdwY7FJ
vRKWph/RoN6O+YmRSK42VlW5HeIdgbA0KsviYQDQZ9jMBrFI0UKFvZ7rAbxeHEhf
ejlRWwunwJRZoNqQtxvYk9vb+grTyDVjp+p0sarj0XZjQ0h0Kk5ONdh2fItqBjV+
TYvLkR0OJ/y/I4SzlHVj3Q==
`protect END_PROTECTED
