`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAE1Yd7kEddb2+YIlSzvqTcs/il7ZC3oeirTlvf4nIIv
Qiw7jUPpaOp7DW3Xc8BHDIARDy5cIwjrGxt/I55AqTloFYPZnEDw8tIq9yWybpa5
jzoM9DS+Q4dMyLfwow3nx1bRMw0CQ0KbvfggCZm23IVrTkb7i/LoDJrvVOSUY1kV
MK0g0PGvvSbsg5u1AibbKa4Jotk9sPilg0qsgHs/L67ASAcYkXcmyJDovdFZJET3
bX16PyR134QhC6H3JDnHVAzbmk4vacIHCuaENLRZzVA/UlffkPJ78jIOhsp3+xwP
/441uxUAoTy7BgL+L7FDcx3SoxRVbVNq4C5/3nO5XeY7z1o0jr/QXBEQVMLndsHg
SqGarPFH65VpeUTaGGjEHK+SgCs5PqhE3APGmdhrjWpTJl0zRv8f3zHR+GYwIk3r
kn08kD0tS99FUGJpc5ZFShBEQsrql5U9zB1p2kE+37zaPLtdpnsybCg/hctmHiE7
`protect END_PROTECTED
