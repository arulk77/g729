`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCiBrR6fijBOakAjjt53UtyGbYjavgrsEbfqEss/tMA2
9OJwpuOdVZCbeR+/ddjPa8OmArltMLifQcmXQjyAkt5PXuyhQ7ySNPC+kmyc8QFA
niIfQ2AsKa8UsTMg1FGWipW4O1zvREPdUhwgmFlO9Nyn+T/UN3phATIudzTx0jJ+
KguQQ+hRyO89A96hK7SugrwDkGRs+1NMI5g4Gl5XJAGfcxNY64d9oDs9/3ZPwmwu
`protect END_PROTECTED
