`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40XWHmKtgiH+642dWjKeyYiGiZf3hxiFhtC5ic1tcU9m
D9QgXy0LUTOBtRKpKczUPqDg7A0KdmjO+Bt9z9mbPZ8N8hC6nRZT9BM8TYso/BSC
y99Q9i8ks87kYizwpZfN+UdRnUWdDEj0I2zGl/ux6nEYCO3yxOQW21wAuXohsafk
VLmoQXf6cFEbyp1oTYw55HWvTNCRneSXR5igDT6bKCoHwkuF8s1wNAQZJhlWmM93
NDgnaxUdmpe6C8UqeUG4eGd5TC9V04TNDGjDZeQ+lnDibznw3RDtvkAaRKoxAOEl
chiTawDC3v8cmHhEZELf3ZfbXGsa4NYGVQixqISNhOTK4Ra3m343X2NoMGR/octz
S6RqyLNUxHEAMvnMgp3nXw==
`protect END_PROTECTED
