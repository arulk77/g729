`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL6RrosO0Bz3l+YezcngZgDCGM03C8mPV+UO2Xuq9/V1
OutuS1sCcnzBpSSCt95XalPPMcs4vrYg858z5z9RUVvzqmQAAwRcM4KyfrchGca3
NJmDP2d8Fgv3HJdIJU1uWEZkOvWx4u2ilo/oqqXV1iDt5f92k25+OgjiJU0dTF7w
8CpzPYSsOjWTPGotKvrd1Hd7XgJ+nWqAUSyab+h5PT97S2EXwUSpwrKLBqK1BxGB
+to94aepJ/pjPKj2JXO8k8d3TcTpfHIwxqXeMvUq7ezoqGCIjcCCx3XPBqujjdOm
FvIexu27+9NyzK3DlannVGb9k18DvpimPWyE3cDZj/5sQVc3ApG1/bI6t0E4VDsR
IsyWHcpGgueKT2yEgrl21XWXwcjFZ5fUaVyQ8g+bwbA82Ojmp797HRrKr1O1zBe5
vHHWXJgD1IbT+jcK4kWwE+NwIna9rt8O9CnRzjhKpLI/KWBk0IgOi1hKhNT9leO2
/DZPSDFhzpth+AAnfQrY70DvnEzpIGA1au61ljn8KJhnOWQPswrW9uYQOVHPQVnu
tz0OtR5kvX4muRSFQx78A6J8jr5cxYKwTwt1GbO5IPqZH7R/QiNksUqKo5mnVEL8
4J7xhjLDdZVSz+R+jFnFWPa4BySqpKsvOIU9ziUMGmonOhLkMCIWCZWWwDdRNLFd
`protect END_PROTECTED
