`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
k58JLsfiwoom55rli2IgVEeuTnDTuAJP+Y8thU7RKF/LavPhvqb31/V2J0q3B1be
ongsr9tQxP3xg3GROEZX/QatYNQeXUz+t3msrS8T/YJxjkBnWAJw6QcwijdRl8Uf
IHrFT4aCKDb6m+sOtcYi+6uyuGZWIAQbx5o+Rt8UeOZkQZgJu6op2bBBY4UivLzk
cvWY0UsOs3JT8MaI5hElpHg8aDcZ0mZqd6eiV/3L4xWefjT/OFctOe71o5LyEOoc
`protect END_PROTECTED
