`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePyZXoq6of6+lgqiv4gT8llvhlik0yoBWozPt4h14caO
w1U/VY9Nr2arSMN7rt1FcNETrbRRwTEC7jM4Ho16CXf19zfBRk7yQKDfHFBuz53h
g6aw1oKlaKTZ/kuMrvZ8wV33B5tOQbw0pDCDwfyhmSkkDUb2G1bE8wNoRKPaZ7R6
83XkBktBmpG57Aw2e4OxyilhbyHNNxMo38HHnyyUYz7d0fvlBVT9JAsPhbPHvidw
/Y7VRiAOMwJJl2GKnm+goU/iS0X3UMDohQJqVupraSrQs2KjA2XS5x0X4qC8rxtu
+JcrTTKWIyi5nv9PFNzwD0lC8W96EejqwAVun24BQ+i4zAYWasNwH23l+RBzIdtO
`protect END_PROTECTED
