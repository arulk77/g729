`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcCFevWkdI9JV97c1eHf9EcQDIqm5XbdXsnd/CDreUo7q
qXs6Vv7mfWzFHmKp3gabjpb4ht3zsu+t3HlYZCJP0c5ZSTV0pMRJhtSUjh9HCmb6
O855djHfPDw7i2s6npmC8wfHHemjwLzk9m0t4btaevFbWHgOXcAEefmD1faBzkrK
2qjh1VT5h3gvhZvKPpPIt2PoD18oqy2n09hkz9N0WIQKgWg6UfQnNUvZivGIqMFz
iYhCa3yMYAQmrzVWGV24FlxNidmkvaI8RNSkiCB3YMQMcQZ93wmE6U9gypA9zEOC
`protect END_PROTECTED
