`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAR1WlUJOpMW1lQCr6Bqop6DHxhNtcZ/EnPKJE4DxGEx1
bwYE7D4I+r1okfG//TXSNraDr0oeYV7fGRl/iBiX8uqJ7J4gQ6vl8pSFNHXpwR50
qnbT8TiRxfwS7+DpRbVqGUYD5ISqNsUUvigQIn2pflwTEThxzg2C+Ft6X7e5RUx0
LKNKc3seDUrmKiFRtlGNN6JnBBaQIxHzt5yR4ebpdoMjFOQ6UJzWKsUMlcuLl8JI
dhh2gZr8imjz2xAiLf9rofa4DPiU2qdjLK/OKtFTipJ0w/UvjwG6MwZyHNPviZ4O
bsmGcg0X2lPmsd84IbCwPQPILZbZBnNjjclEU5BPfAlk1E5ujhu1SE08WddiUXrT
ZyFaJz6N6f8944o0kaJ3yqtFwRzo5aEAMpbXhDunjV81nGa64A74iBUVLlU4EO/C
WiheX9+3R3tT2vzSXfc1+0CW+PZhbHJdCFAhR3wDM7Z4kkvn1rmY/3JnUKgTQjY0
pamVHkn1ORIru5athv1hNscfcU92eG4FxN50HRtT+VtkEoUMy3N2O65ONGvq5aQs
QnHWrjxkNfnzSFLfhhuDWKyWxhMzLLIYg+Zkg8S9IJblJ1f7PCJI/rw0sJDmNaCR
ov3c3eiwL44Zz+5jDssiRU0WCKEbbidV42rMOhGkso6CBnQI93ap+29iIZbOJrsG
cns0XhcnkQY0Fkl0tuAxCg8liEzXroI9n+0SJZd3IpmzOwng4xpIKC0Jxu4LRfW6
H9B1HLCXwttPF4o5zBpC9FAPhxmZNOoHlH5Gu07dkjsReLEGK5X19KPfNs+g7KVs
qL3Qk8Kub4/RdGkpEycjNsmOeiGzXmGHt3AaCcA3J9AsyviDbvBUFk/kvFYYcU8q
8IAsqbMmVIu/zcDCrzLAPeg08f1CZ1wSvC6S+2fprvDVLRAwszf8cv3pNsrH7L9s
jF82RuSWpEP7yozpDqRAal/xyWSafja/WtT871XsZqmX0ZANv1wDbcHX7OWqu2mE
FserOtYZtOFjrdTX+eXOdv2gP1H2gPLJptldUFTGWNOt3bjcJu7G930/HEG45b1n
esmmkIAKop4CnM0jtEEO3UHI1qLi08SSiJF7UGHVfm6yBddJOIPh5iJ1x9P7Iiyi
skwCkTe4gzzuY1D1Cy5nCgvN1lzvbsTItxD8hYg2wgRPUIE+bCoK7p7sKEVPsAAF
aNkSYmY1OH5TTVduU7RBucV6AEcQSf/skDi0baVXNji3GcjWcCqYAQTLdy1ZVuQ0
AAw6QCE2/nZSRutlmHD9ZL66ajqNrS9bf8owvQb/Qs1LZhXS0sGabHD0Hk25SHnu
0I71LbOojA6JX+O069SASibz3PIPpPFNNgA9WevQLojCio2aJwNglcArQt3KVqgD
ONNKZr/T1CrsOXYRX6vZ54yPuXM9byM3cA20nTLBDAx3WdOMbPJYC9jyj6vuCyXx
DQ3ktyFJl6ArKfYhvAkYRx/OT8jytFgbEjKCnWuoe0mbkVSSUKyoMVZaBU8CV9wQ
Z8Plm73IWnuTSW9OWL7DLJvu1V+cbXpokl0NIW8Zq4MFfVi6byV1LS3ZChqjcKNv
bD9FbaVxpysVAw2ymkxdFDowvsKUBddPObBXhVnKb7Tv9J9hQIb+E8vuAoUBT9ws
550oyr8V/4HDkVFqha+j07jDI0gR64NeawlxSXUfBWAAWx8ZgkSeYjXLgW0k6IFE
92ZCLOdDOCWOsue9e1Btj065y8nkfT8/wGkt+YL8LkwUoHNmwVlrssHEkOvLHb33
fb4mEW7KjiIw1MSQZ72hfLwxD+JXoLiFwj3pZxAPJIP8PcLjMaSe96vSO0bSSFgC
NJPtZmF4XHPQFJ+7AMgI3OtQ0wfQXlqCpUWgunMeq/pTj95++sPkNJ4Ulu7rTab1
6EQiGYjY8AhcVRHwS5ErYlZy2Bv6Z/fCfZHJ7kP2quhdKjDXIsPB8CB6Rnsgj235
0z8czSnNFnBOa5d7fJ4Zc1MtP4z7rnQpTvdQluEMHHuKNdyEtctKLPqJVl0I9YK+
glAG+37Ifqn35uFm4qttkX68285j/J5qdeh2w71Cl6FA0qlYjiWD91fTN5KbjmqM
Zb5x3NNAQ40EUsGVXA/OCykmwfniebFuu7d8alAz+7TF4OHvi5vCpsnqvAUKsevc
3lapWlx1tRzMhT4pugVow20d9gc96aFR6EIMx+MNpjML9UIgAmLMGanvkDNos6oe
aN8X5yKHq66ezjSY/LGbBGkXCwVqGsIWjjaQtSJLWe/hW1kAyrRYGLc2tB2HtNbH
PMPaFtIWLwJvZ6aJXguVEa76BCEp314OVMsSN61ASIwrVuiwH1sOJ9LWp3VaAVgP
m0/CamXzScUdUrpzhDtl9502Lsa00uQBoW7Vsh8vt17xsj5La/n3M8PGExcpuPpK
ZjWCf6er0mrMqeffP1CVyw4GJipFe6qmxTTXcVApIfEVFNPedOl0iNtJ19qV6Zvo
0s1vE914heyupHWp1RrcZba2hq4dV8rx+EQ2HeW3rGd8DHJ1lu4F3ulbQ0A5xFUz
rS43/YymnyIi1K/HAGLSs0xTWSiHAMKIpGX+O/+116DbvbgBN6W9bEvNscoE+JB0
IL/d3d6hXJ1tHAiPrQ6W0J1GG06DrCCffLGsyCAawVBYHtB31Covz4k3YgHwyGHA
OfPJX/XlDUTGTO0oj4nJUeoaBgMwUJeJzoyIVUhsXU7fIsLZimRoU0a2AQjVdtst
7MHzvcdf/jdznOJBobIPFi8giYyRJVlN0t3f2Y8aARUqb/WDuKeBjOjFzhhOdxI7
`protect END_PROTECTED
