`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aXUzADGnWK/r+1zAMKCamwxUD3e7Bvhe3nJOi2L9BueVsF5DHhbU2Yf34wGmR63I
/OCiwFcEPiZMGpagLVbMGBVr88JOw2jNNLfikArEdddUYzG5AkVHSwXRTviCwgh/
`protect END_PROTECTED
