`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xi1qicUzXiyW1keCI/U0Xa+pkHuv2ZIWoSPsjy5WcdB
glE8NntI4E7yCRSHuE7eVs1u/8eM6YKHi9zdxywGx6jsenZADQBHJgS+qzN8aKQ+
qo8TAI4m4YyrWJYm6ranGXuTlMAS+nQYw2SGvCRfMVv3ZFvWHYlTyoFBdqPUP9A/
V8pA6RLVQd6Bng+ewZ6axWmhdRF1MVjNeWthZ2wrwlzX7/Mw27Maw/Dz0r1O2Xuc
kGP2o31Pjvtt05q2vvovZwIA+5OZnaXElW1GKoj0l1hxrfyKibAzVTyophgaJKRi
83zAcZyvQhwphN7SQ/YTzw==
`protect END_PROTECTED
