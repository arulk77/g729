`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGvPzHSFIAAoU+t19J+EZ3PgveTUaQqWuOAQzTyeiY80
obhHiYW8813WZvKKWZOTb963aaRoG1SGNBFLDfUQq9y9XiKSaRt5Njsx1E4SGwIf
/ZqNmmTwzHs5jdfVUfekjdy//TPIXyJk5fI8JVmOHNF8BwLWECZeZrHCuvlMtNez
cggMniK0CAm/Un6wE31yspxFfcd/3zIsLGoDG8P9/1xcn0cANc2sCMLL2s3HUz4o
U2Y/6brQ+4NkAm9lypafckbOZyeBpPbw6dLwzC+DTQjiv95zelX1EDnn/udA78AC
Zda4mzQUxy473s09XzlRFrWZWTWU0xYxpWzSYnEtbdF/YlvTijWbHrpSeOBBzapz
BIdyPtYkfsP7DYikHr9khvzPL6R/owMsExZzjIVA5jybkQNDoPsVYTkU7BknVz/S
V4q2+qEQRdnQGGq4rCSxXZf7or87n7OZxlrtHXHoGDF8N9qDSX61U2itohu5iHND
`protect END_PROTECTED
