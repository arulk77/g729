`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lCoCthqxC3Eq5TaEgjoIsV2/3mhbhLGFhYQm1oOwoAJ7V3z88pR0KP3Hb/q7UZyM
RzRIx+v4r9YvwE7K0KYD8HImI7sOBT4BMi4DquiuqBAJLc4tpmNMeEAvWwAxPbmn
8tgtEO+16c0xAv6IHlR3BtycKjQwCL1xcLUVVT0U+Qg=
`protect END_PROTECTED
