`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu449DSPHrOvVgYWwvCVu8QalmHWtCQJ4xnAIpT7jcF0yd
5giE/iX4OfpzeR2TSFzAqLJlw6WRJSniMvn4jp3Qo3iIeQbF2FgEmRiKmLOVM8ij
VLrpGwYrnEN+/gUyjmirEjMciI1ttwUGSSDLUKIbRmUHQvcREkuhaK+FAIkVeqra
azOhbX9v/F4CcPbL8UUZueh2m0H8FnVOXNlCFPwGtmTy5q33oYYAObgXa2PDpZED
oKZhvAO7N2y+Hp+TTkUqcpQRTe8ax0NA7GTdlYN3RtNFaymreQF5rnaa3sCLyJLz
3iSKHSo1CEjHDmLsJ5ukQg==
`protect END_PROTECTED
