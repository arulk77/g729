`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMfgjAyT1MTPCgCfyeQcmxz9rxHjEid+M3Miqw7W/xNG
mz0xy9cp5V9S9rZRZ4McVqJBd6SVPp765yCWL+uWDEowh6k9qtujCxS/MzvY/x6Q
xBrujCUXDO6Xhw5Ao/DmAR3FkPb2dfGWNvtRSmNo7CSxRFhIgN0Bo8p3dfCRaOB7
h7jyHVLRiP9f4eplockfwPmO45tEi1LPt1/gXOZVtHr9PbKMUAJ6Q4y9XUY+8sh/
aeP288167hvYcBjMjXhE2Gr+hRvmilg4F1xjeHUWnTZhXCgg5jH9EqBiCf7Y1xNX
+2rdGO3LsguWWIZWPtVsduM6DfE4SJpMEGQhQb7GF/maeGbeRqlSakKdYG+03nER
0a0x3R3il28gVZ/1fetPE57fEeSiiiDldKptJatAFVXCI/YWuSqD45hA30HDiZBI
nX4DZvLS2RU0yMlHIOaG99khklYlpwmurAKdtWEGEDJZ/UYyDLieeYuYDWq4MymZ
v+CWga00cQKHu8ahYJ6pgrp1RNFvzY8MNhN/7ODGfHfolBlRa5hPmqGSTdnCGoh5
9H3dIUKBsc1nZFtRE/BdM/hpqe95EO2FtdTc6c6H+xGjO1148/UoqTbqq8ccDClv
lFN3r3dCjih3wuNg5o/F4NubtDGfuu4ygzJ9ruTz+rFuGWtGd8l5Vy65DCqfFAlT
BHi7Swsghc1fyk3fBH8OMeSnRUz061qLs+G54yBETiTcl2Maj7jmyBSiClabeH8d
uMm+HdtVm88vQDgKDByEbedFIfyK7lr5YtCrP3PvCEPdudRO0hsSoLzJTePNJjpc
4HX6Q2fUubH3Jo46aJ9ayo9FgCo7tgzadE+8kl8Zgb8=
`protect END_PROTECTED
