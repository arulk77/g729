`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1HXC+aLVpXZ0dZT4W++R47owIPO3sPXct65OBv3sCgtx3KNsViWdCyLNRJeH5WCR
Har/6I1XwQA/0twuqofLAJ329onIgnGfmQBGIf/JdIr4j62mbmesUBzpgq6oke81
GLos5lJ3GDDSgrm9mAH4u5oA1RTOTnD+02aGfxOfXFd49D1Z4cb4kHxyIHmrjXm1
emwR5th0Zo2lZtiDt7xP74+d0wihl0G9MQbySl3W8sjLuTF0Paf9HGqypthN5Hru
H4YE1pxbLpnxksgUUpSSCMbaVS9HJvEwns4DVH1hLOZlgYASubL4jr/fGkYvjhXP
usk1bGnS11Fu2x7hgBfg7MDahChZKXyh4uVgwizr8IuIymEpkKcoXeQ6ig7AGITq
3xYRBEsj0mK3wClDy/vw8E7+lpTQF1TIllkGdXif8OtQeiojpEmCmF7RiknAN/xO
XOatDpNw6rGPTX9ZvQ4o7H6HDcAaiHV9o/8Yqp21W0+k/g2phnNQug8GSX2MfbDs
iJpd284D7qCH6mZ3VkWa0jHonRDW/7eLphQbfFaQDnvQ5PJ4hKUpkj2b4Ox+3ixi
WtgY18CKBqUXUogO5t/Sn7n8vNAdrfJ9i7oHX7PrybU7AaTO3ZYaE0YEtDAChNJ1
s78c0hPPJNUvIG3jD6L7HMhyWka/pEBlBEa0lrXUKXPTGhRgzEYaXb5k+jy4ty3V
ti1VhcYKkomBuAFpR/MwIQ==
`protect END_PROTECTED
