`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL89bFREAXvPjIM+3hgDrwX5DodcgWMEuAAEdTfUJQ06/Q
snEyqTyOXk66xy2R56KB2z7qUYYbNZOzTUlY7qoch0dyiDNrHHAmcrP7MMtZiQ3l
cu0/yxqobhfUU0KChYooMlnNqQJMoF8flGTGfTNyL42aveG+FrdkGvMQSut+R5wz
2s4UmLM3ZmiwyAmYmBsnS6OU0KMQ2r8Uox3AQw1MATg=
`protect END_PROTECTED
