`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePV0a7Aj/RRHNxrDHNuGSgXYEXWq2MRt78+CCLYjZifF
ey4CET+WY5oTzB0D1Wsa07lcs9Zp0mmnjguUvEjeQ/ZC30Hf2QVmFYUqp3Csuiyp
KUl6NlB3ZIVPRUROxt3K8CV7INQioH8vS5nuXvOHV2ZXHIC/PnMQCy3QYXYs9Lfi
kISnnkM9s6BOw/07B+Day9iArhyy00juHlzZ/HXL6vjf3b06QT0Ox5YUCw6LSoQq
vEjE8jyz+m3SekkljXScNaC4F7Ml9HLmE/YYxUo6SAbi2ZXdiom8pnWjPEfLxtCD
Drz+ASLYzbCqkZv6wuO1wCHRYpSFB5OWJ3dAmQs8SCi+6d199yI3VSPT4x7b9bf/
FbBLAIfxZ1r6Ywrgi+VEKxhCXMuek2lmL6gNa/LhuhYclpFTNIh8bipoaFBecZ5L
zE4CH3CoxMro+mwm+BTE6/9n/jj+f7psV5d9RmheVmrmVRmz9pEzF1P7R3CihanU
AjMzZen/XT9WiIXIx1/2lw==
`protect END_PROTECTED
