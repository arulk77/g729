`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C7DyvuW7Rxjej+ZAI7e2qDLb7yK9cDYBxEIe8Vw9DQGu
kn9nQmv3/1W2SOVvJ7p0jkmV8469rXtPtL9JP1FLAstl18MT6zDA2L2gitNPGvEc
zqJOC8MbtLF45yQyIaRjehNslDml5O5adlN7BsNsCHK8saB6D2yQF7mJtxpoB1E+
9ecbijjBRTrGcKIycup0zI0R5jZM+27Ym8MSIu4DFbQlGzyu9sQqzF28PYSzOd47
Jgnuo3mrhv07YDBhbU3PZ9dFkDwpYg40PE52Q+f4ySZnGsSYG3GRVnpszh1hAqdH
wCJ5JUD9Fe+4rmqvhaxVxC9Mmm0qCR58zg02Dhn2xKl17q10MuH0nZPqcwgiQG+m
Lyq671eUetPdxVpYPjvO1gV/YAcOMB4eGQF1LqVHajRk0CufXP4ixmOiiwM8xld3
PpFIkz9V4OR/20KCn21pZYDVTgazRcFI58s+xDEwCX+QJjLn7K2BCMwEPUpDa8Ow
Ylm2ntydNOVxLyasKk4/vy9UOJ5OoJkmtZXNhKSuxL5OBy705Y8ynJU5zUNwjch3
TvZ4Nu14T4+cf4DjOAsJg3ZAs38l6RU0u/gjnvVaPEsEyBpBLmTvV/fU3p2oFNTK
WY3Vv7KBZAt0bg6QGNYsaV/ezKi64MQcFn31FIpvECQytQsvRhQmAt50BmOGYzuD
a0eWgOCok5ddaz+ba3xKYU/E0++KCHKi214aYPfse0iLWJw9ccCUtQqt+9MH7+0B
mD5VF+B1f6LW92II0IvvvAEfdJWInBRTrTprSdNrnbMHJ/jwFthutgLy7/q67/Eo
wqymMUf7yX4W5RyH/kzYNYhieygu10p+2TKQDjwGXmjm7inR7QcaqB/i1Co2vASx
u9LiKsbL6/Cc/QDG8VSWIxj2OzmygPTEtnalGBWTBfDrF+FVLlYVUKZvMofbpAV3
rRfAX2nD4HDMqFCexEO9ECRjuPbQJSyOg9bQDHSeRaNCN/Sr8UGapX/pAenahdi6
+kpDpOj2m4SdB82//D+MTsJP074du4UzE0IbYY6uwBp40oxD2NydpEXwqGOJGufg
wEQFbkUN+WRZgUGgZg/3Orv8TfpPcABTKxm2N70be94eNbuzO5tnj4tk1hZt+lnf
c2I+B7jLAlh1rohoXAvUUJiEIbSOL8GAZBSDDOoaj8Az42wi1PKn4QieycwxYq+H
dTRaHnyzGdI1dl0e9j4XPjiHkKL9QBxiEhkWjmLgzBbCEy6Q1K765ckUpLx5tKpZ
9KAkMza5Vw6FiK0lWPA2pdO85+R0quS4lAIXmN9fXsj/eaEvtlsuTptsBKWy2/jC
5EEeWKNbOpvavNQ/TEGHgsk9x/FDxxAi+PIFZzdddPQSGSkxPN132b8OHCiENWah
5yP3P8JECN93XL2ZxB90jB6YabdJFKP1UbYLHyy0bguU+qYUqWlfEGbz1xr3geRp
l7scwjpvnnhfGUuWa0hNWQJ7dqYPne3PpntP0FSwV2JsaK8+j7CbYE/j5bkQz9Yq
HU7fmWIufLPyoQsLJB4Lm68KyyeAsXh3UHETu67dCnCHANVkBdBsc7zCIeoFwtGH
GiNFY4HzhHIlPZ5K9/5kla41RlPI810dXdKScVMCnrS6Zrr4XWLNjT7afH4JDjWz
AsTileqF4sXSnWPxtiahJ3jSqaCZchTfJVDjINaw40NFDCQvGtHcsysFn1tD8NZK
Lt/WT267Ep+/YgQ8qMceX4kurXYDPavxv9MS1dS/sMg5B1QG/Q25qlMy5ZZpAko0
6PYu+aHSH6pQxWbi4zlAVx1B6A3BrqRbf3gLUDSCSVMQb0rIf2tYbSF5zajmbwMq
7M/GOrKszVKs1r5bpih0XLN8ZR/3MrfDDjtAgsfpJAuOFg6mED3c27zGXLpGk7yp
OolLnWG7S1kYVm2i2evjMjwapy5i3wj6aQGjJfI1SkiK/qT06QmUVQo6Fw7lyYjm
FbkEgyzBTXwN5yZVo7is3n1CcnHjrStoHyqKcmy1KY2YkF6P0s3LMVwepNtaZldK
mdVa/tNQLVoLjxrDbghUTHREjivk5k4MGnP8iAcs76o9vhQN0qByrCIgns44TMxo
O0+FqddhNbLJX1OS1Zpg+b8vu+Yjxo09oPtJ+9d4dNvDklvm1KD9CA/2NuGd4zXp
8NHh6g8rc7CiJIeZbZ1/edIuH/ePJOWITgyrB7WRcPX8NdqcpFaOh/vGabBp/x+A
yqYV/AhfQnQOKfQS/5iIzf1c2kJMsLhAz2gjsAb0HHH3mv+otugVPf2Bh54hbaMn
0Xk+fgpoh4qWAKkpNJAXPs50QYGAQ4Y6K2qPK2X0Wl3cnaoUqAc5z29VDllbPwGN
Op2s6lEw68xYZr+NlUyoHaISvEiRINHyhg7l9svbICX+UJ0nUuY8DF1BVllmZ+zp
q8yTvxAfY9qd5CNH1twrnZVSZFYZYJwfwcYNL79ieFLX5dmWFZw/1gPTEurfGImE
fq3kBF/AMHXaLFWolZHZyoHoxHOIpf2rfVeobnnnin1U/CnoNZ4nux7W1k417IzL
j/+cM9hJ7TUIL5o5YFq46SUXflnzRkMDQauiLF/menfWK2EKh80sV3aZYU/fw3rR
ehageHHTtCvsWyuhI6ktdcq7FSd1lOsRHe1O0PGBRVXim/jeouEBsiHIhXswcECP
VocFGNDU2fBZr6uupH8aclYkvzpfUvPnZJXXD0HGm1AGjKeLhL5fNakE/ApUfCk/
LthLko0PHfCo2XAq8kktnw==
`protect END_PROTECTED
