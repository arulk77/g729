`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL83TFqqM5JZf1WEt2arccWJfC8CDGnodwH2pC3oM8NVIC
uf+jaaLepN6RIErX320aTZYjEhlD0xuUhYiMVtOYbDnZHuDQQCxqrotjdvFcqEYr
mY/RnYjmFu3+joOSA4ocfRBzDcU+9R3WWKquk0bjH1o2drfu8fwZeUXSxooQFyxA
Ui8IWoSDomEJ6DjdtRMLhPiY7k6Ol2iAQ8Ovv3I054glahxUUbqxZ7eWn4oj89PD
nTBAfuw7ih98x4zeXeWa5RspoSqE8OMdcIKqgjrUYQeO7F/j7gIrV5XYJRLHz+SZ
uWoVuhTZe1ASC3wNHjACoKc6waHROaIHz0JzhQJe+uU4AzdUQLHsfE6BKI4N38nM
vg3MPM5eqQTS6Tyv322xccQ+sAvG0ZicpXy+U85t/JGC0FQN8IhcFL+HIsF7OsoK
qDnssqOvpGjCq5nau2GSpocE7mh5mpZ3VgOZuBHVja8BPxICVLJ1OYV8U2p3OiOe
5LSKu3a3Rxz4lvpzT18R3xZeJwL63fWDJIKfWGq/qmInH6b+fagqxcVpN3MK0ZwW
3bm7hlr5X+Pa+toqGnC/PKqPi9NbAwjPyXZHo5TrubXtl9Kv+0+qj4NLXP5FOU6u
DZoHcSHIm/ol16y5wfvtsegA0ZO2Sq1rmZzafOPbVfRD/KF3oJ+T8Tzav86iDE6x
wJqi1AD5t5ZwPLBWlxWa6/6+rr9OjctkUQqmI3VOSUoz1e/1iMyD2FNNl5LIZH+U
dD7t4+jJY32L2PD8A8j1Uu7jyPuJ8SVQGVu66t3P4nhbcGhqrH4XeLfDM2MVLQsd
U+UGkfOsnPfBBCOs1bDUc9erThZdsI+2JhmE1j5Q6LztqtUE/4pjAMYGF+nNm2Fz
V54CM9OVJVUyDNWhnxodJuAXHVUB/Femp6MJxiUmm+JmwSn5TvEeIJjJztkkr43h
axk/N7ZRH/B29DPKIaP0BGqWbTIoJS3faWj25/qZz62UIrx4ZOCtldTQiaX2kGE3
rWE+QMAkYrqbXfJyfezJK2JCUNd62yljy3/BPJ+nz27KnMQXajH/GYLpEvP+CwSy
HcGn8oXlv35Tpl1/Ccef2cyS5DDHg83/3muUX6fGSnbD0sR3WXWLLuZM8eHJIcLd
TUkc8yEkdF7xrWExVZTcIv9I8cuomWGIvrqZXlCqsw/uHj4SmWjgHftMFQ7IdYIH
jcHKdo8gYS3mGtiZMijz6MmRlu6B+nBPs52QuQZm9is6mnpkduvQiZp+zJPQdlws
A2gEicoDMVN8qV6AyYKN+uSr/8FSw21tXwYJE5LU8jVUyE2OSNxb29oCR2z6zEwk
zTtcMGHC54lSOeQLus6I59NcArojZfq+oKBKTa/8BXUgWtJvA2Pu2iXgYJL5rM1I
sfuPzzo2GUMqAyfcsml898zArbZBe+tpA6rKVthlzqox3i9XI4KBogziMMRhTTvZ
469G/UwVbIs8hAIsyzaE8QKYEtQ7i05X5mer+JMcrIl18Dy14qnqCSi+NT3LcIc1
WU72BzitN5tWnhfKtTwHa39z23nxP5g8AXLWhUlOBLHkSvWdtp8UTHedOUDTmjeu
11v7YY2q1w1YUGR/cqjWIXKuz5m4odQtqDIoi6cJ28GexvHieoMj8H/qGI88ZRPt
RnGoaLHBf6kgQgreXN+0QlIRYjxKUz8df4f4n8tuC4ToOjfhGKkNaXYoHc1cDnrr
0X1yOwdFW1O/5FKXz3FSACA2iDTy5ss7tbfW5JwfWmCxq2PEI0vcBPZ78IQJsFO6
MQa8TitkGX/7Mzts8HQnaOQVs/LNzgyjmycENEzUiEzT5YiEAvzzF+SPvWGc77Gk
m03GAqhmNOddZHclbWBz5tpCVhWSWFbKhlzesniOLGwruptRWPCmuS0MiR077rrZ
YgDeaVom3rAm/vFZ9rmKTNheW4xWovw8xA+dqbAIuorY6ge9XGWAhDi/+wjl2JKo
MVez9xJ5qfVkKL9IKXMhEAaVf9W9f/1EX7YysL9aci9NpywITjQZLdaLvw5y19Q7
ni8B5LbpIR9ry7rc7udWn3E+Jw35tNs7+anzcu/GIynN79srUSMFm07orFiW1qmU
/tiiex0NY2ktYzba9r7A2X9Ds2nBo7PQuKcZO9lf5AVvWZ82H7OMVN/58fiLz9c9
hMFCxsyJ5q0M8qQNjTpJH5d7uL5t5P5ZuPxma8ji5UsABiq9j7BuSSkN5MzvPQAg
dKA2rE/TC6/GmCrycvmq3DtKU8UFOESij65MwtlrnyYA2DhbXXd7VyP0t6zyptQF
JvfO+cI1ZXtFc5egvNfw9uXn3PQtBWEZ1G0BIVlwN2BFPJXiRcm8XmJB1vz85S1n
Q+OC/ybgFhq2EJNBszmjNrpHK7fxfOGB6+g3Zj5y8V2UfR2VZh8HPUNQVGMp5nQe
QJ5xKG/2zbDS+rP3vT5MR/r4gQKdqKqa8UA3vY1+q4u2uIWidmfxNlVEuTbKmRhR
BT2tVt0ibdMLfxNpJxe4B67AcaDlWhmSN5iuSqTl6b4XxbXNwm3NvP9kgRMKfEV/
jIQHoA7j9JH5s2wj3DdUaM09HBAzJiI5EQpWuzGBh3yLI/VPhcym7qpH4AYi3iE2
9h0NSfdo3iQqd4F3Vd68VuoHBXCHrgDWdVbCFsej9nT0cjTJHrdOOsR6jOjdIrJu
RDE6AFoqKk/4pB+T9cWmsQZbr/Si5m9p67DT5O3BDRh249mMGLwiyqQRcBr3gygv
gs/xmXsluFO+MWP1syp/YPjjkjaSOVpjktIWS/kjW1k7omuNUusQtoxfdS7Uo4mn
/BtQs8D+JkxdPVOcw7T+MyAsUXKQKT2SkM6W8+AbSxb9QxdGSRnTqyEbUCNiwdAM
5K/t302PIzinmK7amjKVVFxRG7jNkXSM7VSZQ0jibaTQ+85vGk7Q9XrIASXThFjR
kt4YwHYxjJ2eF5TLHBr7VhTBD+ir7CsGzEq17AWy1zYshCALKWy744Rn50/qTJIS
empA1exIe61OyateAZEScmLoZYBYsoVJug6rDaVpFBked19ivCNt0pPHOKiorrid
JuO66RNhvKitnRoZDpO5NrZPEuEPVrjG1SzhXHhM9SR0WwOvIrq2mKkremb70Qmb
RUqErvT6TCW6XWdzzcqG/AmwlxwgHj+Jn6xN76x+pKoIqU+Aa7o5PXAMRUgHnCkA
SolKHT0Nvw9olFPvecmH7KUWTgnmyVlaxclCgQvSRQY0QVMLJ94O9cxl+w/+J3kQ
/KtCNhwiWaFmslUkEUMJvc1lZ8QmpvDVEWGrvQ9UWfVicRlW74APXSYNmv1gDRkj
QlXGz04X36fGgB+Cgo6kZclU1RA/bgq+joov7F7Uc/m12b1QiLMcXPBtyk8w2I2Y
PdQaewN2at+03S3XnjOjenV0S8Np/+tGqabWhDV1k17v2a3vW8h9QZ4fXDta+fR7
Ck6e2IKPD8nCNhr1oazaz1jLdhPoKFvig+aYTxeuYVxkKJI+YCfAaJKbQwoJUPvI
H3QB5coRXY/Dk925Kbu2r8j+k7P1MWe4iNsRjDeHWiMrDLefDyFrrNXdozGe+vtj
0W27miuheOMCBMu0Q0N307ygoceiUcAjVgtZiVkvm+U=
`protect END_PROTECTED
