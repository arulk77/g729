`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49++5+C1IAr0C2P1/ZTH5MUKzjlXCu/a9h3zRepZlFEv
3U9ksEFHZ/bHlip2TiXrZj6vkLsx+EP4RQxwo9Aqr4sS+wrsun4d+nkdQkWYI7fn
388uNoawrBSR5pgcQgvVnAgPTOwONeDKjvPMNUSWQSQFlnvEj3VPQy0pTxzv+e5m
z3UT/E+Ybv9cY1z/lfhL1V8M+4yBx4tEJL3NEvZWsElmD5xS87J7gcqojDPly4Pv
1huuX+Dm+VermXbolqkxVBBo2EcEY8SSq8aBOe6CX4g=
`protect END_PROTECTED
