`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45l1aWjAIOVqfoq5e7Ndt1884iLrDlN9nyJgHbltMGgb
uPU5ll6T4/Hh43fqPgsV8rcMV+CYzMJMX21KHnTlL/Hy3J+zLwxWhmhtgfYA1pc9
Sis2aGtDAaNQTCF0JL9teTwul+74HPwJruh7fzSOiJOE+FnZ1UGMR0uufFEsOhKJ
j/0WMnq+YgY7zEi9QU/kOx+al2BSYR9YPo3WrOxAf0ux+unsBFH/qEUDDrM/CP7u
e1B8yADILTLB6DUMVxuNKIpsz0SsuJy0bfhRNWU8But+RouYVHQVnf2reuEjrdRD
8d9ZKVA9GMtyaL9NHfRNf3FeunVaQyE3qiBRkka4eyI1itwv+rCIFRGFZMk+2MJe
XZr88q1C7nLFgs2XTBvPJQ==
`protect END_PROTECTED
