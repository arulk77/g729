`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBTGWTHB/D2MhOY6BeO+0Wj0uRe8d9cQeNvSe3kTJbTW
BHi6K+aQLRcZXsZfjsMnmev3AaFNwpaIyqN0ySukuJhipDcGawsSGiyFT/76MoB/
aGn8CN6wpqftShNAZ9P4tTdYIA+qI0+n7jSy1WBckQgu7KhZToKblUr4ZGnccpEt
GlN4h58JDCt80fhjJkVC1IXYz4uCG0eTeLFyaArPit8IVF2sQ+sf37t9ktJRnvrK
`protect END_PROTECTED
