`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFCU/HKtD4mzuG9TvMpZzq2fDRIWIJ2TeSpmA5I/kL1l
KJwGC0HJ0rweLj2RYqrxK6l3a5oUEvA3IW8POsZA36u3rMJT8rY2DukPl8utTtXQ
G3Vjj7aTZo840zp01/lTI4XErL1MA1CoXmEd20rBoebGofAf6ZwQGW/ReAjyLp3J
+qoesmZw66U82bWjNQf/AKnxbXLt4LtpLjUXUsudWVg+ChCsCClakyHUNfrWAopy
f+q8C/Msdc/OX4ZP/nG2+TxSukLxpAaKOX2Q8OrhWShwlDlIHR1iaTdqwIHye2/x
sd0kZgJX19GWREVUo0IvXOIOKsWRaGT/ujfz+2fjTRihSZZ08qYnAQVSFyItdL/8
Rjt8u/BmPZV0g9aceGfrUk7TYRUTNXKDy1GyKZxrGDRUUmNEmdcCJzZiOe6Jaaiu
cYzjOAj+ZMEhgj0AgFzilC4BxkqG86Pdrfn/GYV5E09s371/ugrv5uNq5mJlji8v
`protect END_PROTECTED
