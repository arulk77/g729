`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RH3cFFctB4WP0QKOIk74frd/15DoLoS7uz8JdpuD4l7oCitBy5VAD0lNP5wGZ2s4
lZKWgAutZzolzW5YsWQ4h7GdF8hGT3SQ8KLF35VWHoWkNfIji7EICCxMgEiJ+2YY
tFl8qnZtoixUtmfnWJ+d8cUqMGO5tloKlxL8NNa32tjAVsRGbncqF0zgkkzg1RbK
FgY4O2X/XoOBSBIWCXnjqtVibI80U9MfL3SdjqcKIMU2YJkSHbmEhgsYIbEkNI2R
qECm6MGaOC1/geokO11F0CR7a4amfcb2bKdPIQEPvRAAWA5gbKyv3t9fsXLlzf75
DYX1MWMf1bRHEvxvmu04WMr4+22fEx0ODldwteSJOMLxN2AFsvT0Q/JtCYoUBreG
zOlJa5JtpwI4cK+S9WAojPJX7dAUVyb/qD3VhzZVTnI=
`protect END_PROTECTED
