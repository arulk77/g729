`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEjie+IQ62GRkgOum00ojfvfkm3ssjZpaIu7YpvWqmuR
ty28C63Bn1Z09TEbLrFfM9xas3H/8sW9EAW5qKSO6JOu1udoWKdXlMUPVQ6QzIYo
BCxRe3POTDHuI/4+LWnBbuQyyDSYWc3XS1QsbVEOUYSuHbDQazRhPP3u8vcHBHyC
h49MXt8GuGDcgX5drl68rA==
`protect END_PROTECTED
