`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDdIzJQWzUj//z9yD+q3Iw9z4dOkB3JKoZWCHnyEKeFD
5X+H2l+fsQ9qc4tjU7QaEw2C12GagggR2XfypxNpMq0//lC83dpQlzIQAAflIi1j
rzE50zzjpwtWIM20cMZrvUnMf8ckysokcxx49x5sEJQ/qk+krxGYYLaHKomYEKgj
c78KoNeOPAIZrfjZ6ZbY3aJsLe0gv2DLXHiuGyViNXX85B3t+07hSbiL7xsX6y0M
XRixS7PQTMqcjX9OZvH6o61lPZDmskgFy+j85BFC9ArAlskV1+ydvMk3jhn8Bi3h
p0H0Dx7utuHbT3cO3CFaMPRAPqBlvEzxtH+9hY9aFqP2nUea4clAoKuXnh749vjC
AVLvNrOUqz59X9bC6+f9X2BYplzrsODs/DB2RzPo2Kl0TBHf5GkY8PH2vdlgWiN2
MPvt1wCTd29kKvr/BebMAyfM1hXkVPmazcVDrTEe5IUuFymtRRUePrqAw9IXjOAu
`protect END_PROTECTED
