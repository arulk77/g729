`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNN4NpVo/x4they2tk6Pl9tf7/PRrKa7QME5skQPk7Ba
fjtBnKNg53KnbvOg1voVBO8jIM1P0g/v50u4csWShwV+e+rJOj9vwu3Wl2xse7lk
B32QPIJ2JJ/zItiWpaspQH7Fk/Txz27QJL4r9DzscE+cutJ1nBwJaqNayWFF9+Cu
G0/CcqlzXpTueZ8EkgzfXsAqQJ5UCwXLJEH/vWauz5PodX+UmAyvoKqkgDdH9vbq
3XnpTBsuHvuYpy2mycMhePxYjPtMsHLk55LuQkP2kIeyoRdaz6UaVjeBzZ1YUicQ
Q6h4ICtGnK+Sgwnui/+BVT0ETXw1z9ki26tcMeQHnyoLkV3HvsGIVl+EaPYiMoxr
aGkQ5uGkj9U8OJ/f3qZbruEXvJCCo07doVnlNEJg83RyZYikHaJXN/YL4lTfOt57
eoCoikeQwkhjwu/YNXkasFDC3+Wib+JKz6njEQLKyM8BMXvy9NZY/9zc2zT4plu6
V7H6cu/NcpfvMX+0fpVQpAZwPnNgggLAdxpyNh3JDu94Zhcq/YJBBbtZsXNNwOBI
wJQJoB/bbzu3WbJlq7P6h/F4zxOfR/dASwuRHqGuVJD5Ueio5akaEhRhR0wG0LW5
rHmsJlKgHNnXQPYXJnnQvnROTI6xD4OAqdeMKOORGF1aN2x/5cRDkas5zP5AepxG
`protect END_PROTECTED
