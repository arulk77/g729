`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIGeyYNJDGKgnJm89uiPR86D/8BCDwYcW4jaVFEtpRnE
/mTji0REnBZ+hG/Z+HZ1nX+H7UkFedmM3gcW+6bM7TF0fGRJ94sIyqFZ0ZUDU2xL
9RcVl23RUcvBJyax95xilG2XH6MZEua5BdMIj6atRbBbg+GEKWLkBJUrNf5+OboJ
sCmZPwcM0EK+WWjudCf85YwHwstP9YRibDJJq4RdGlYUmYZw7GIo5+WILlBY1nyE
RTgQHA/F7ziqxG3eRI2jOzv1xmEPk6fvX9ZhVxRnMMso6ZSwp7YfaY3cAR8cDEsY
8fVK7PNXtSQIvj6jz/rRMSxUPLSd2g4ftrqG5dZZhSHP6YioBICQjr02rUocZDEg
kzW0F/4JV8RexDTCYFXS/IlcUY4JjUxNofrI4LE9Wn3zz659KGJ34rSviEusq81G
JCOT7XYfZMMsb3Wu/HGFbzuaJ3Wd3wDnPpKwwGjWxDqxeUzXFaM5IO0a4q9Xrzyg
kjsmEt2dEuHvLSjCKAbwL+wo0Gb2ctTiKNa7lsuE4yCRTpXARXcbtDdlwGAYzRm7
`protect END_PROTECTED
