`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM0AvUhhpSIFWx2y9INameFGhMl7LGIpIaWXSUWuf8WE
2WOi4PMKwc+4RWw0+P+AY+cEE+oekIc8uR7jNBH9dxUesHAilobqdlsqAoTpfONs
l0jT+g7xVuyCdxDdCaa8s7npAYojGc8vTCKUMNUauFIeOlU82oEGj8Q5Y+irtGN2
aFsFjcDyn0JkMgKlLCVCslXVAK2Mil0o7gvdzdsCIXVKeRr9tbNCtUT+LAEzqd93
OYyRuUjuoCjXWTFdnXjErlbQl4cva/8QwtpiME/G43Mr5NYDSDeb7VVhPImBq76M
yCkwnTM3iry8HDBaEb81/3gg9Oe4syQdZlK1780YNwr6Wow1GFanl9ZyHHvUuuOB
cE1OJpZqZPt6FtBpoibfX8EcdFpWRqyjY5HsxDpLHqWWy3gz8pIqT0YqdHQ6J3LV
suQNvjhYHrFj9fduX5kPks8GYT6ISoSQexBrNaZU3u3Ml2GyqKZMRz+HrVnCw1Do
uSwV4qK0Rl7Iy52xQS0Gu8IspvjnVIJhGqG/dXPYyCezP+BXOGO2+RGCaBwHf7nS
`protect END_PROTECTED
