`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFlJYdLeibNh6Wk3y5GlbUoTinv1TxLK8zL5CKRxrkq4
qiHr/st/GaMs1hO9XsoMI1zfHjJn7s1Tdv6pVr5A7f/sCeLOaEic+EzXJIiWmRiM
cu3aXLXK2nfr75A86SbHKLdZa0buhhQUgZGx4jv+tdizCERF/eVSbv8IkSGda2/1
cHOVt1vAtUj61kQCjytsEpNaRGj8JFQEOKNVlXKSTata91bFOiQo56pun5TGAOOp
PlMMROMRRVk9knp1sY/gZ39ccXyF6hGD+Ur+NFgWCcWH+lTVwrw4osDUANoJX8ym
nBU3xB0nKlmpIHXM12a3LYRDI61YWa6H9D/fcCBeqrmNejOUeejDEqBJv4lC0yKy
lDlXtgBkpSoW8E2OAFE/qhL/WVslHyUN5hGHQHXVF0kDBmJabSVDMkbHHlEH9+19
Y831cwHAMCInV3OlzQbX3vUxSpTNWPZnN+3t9Gvklt3Mn7AgACnrEpBrmhyY2U/x
KEpNzq4yaX2/SVjvcj37wJvhqbIle5EfD669Fct7X7IWIn3jHEA/ygms8RsD9eZ8
/o0OOGZlxFQ/jJw8nOrlPJeOjr8gVWgH8fUWTqhGNX5w/E2cYgmhrIonem+GILyB
2bTRa3iIGcxenhLxzjdhIRpIOUoNaRGMfE+DZy11xmOJp5csU0qjo7rWCF4rLft0
lYv43GZeXGkRrkCdrj905mciWS6agJCGI8f4oMRUaeQznAQ75J0eJi1616ypOugL
XB4ffm09lBpklrMNNkuMHH+yfAr8FfKT6ojav/6VoBOuzvegvkDzeVIm3Ilyhls7
SXtTdIrniXWTczXALoX1xQ==
`protect END_PROTECTED
