`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NlMCMefCUkLXs5xCDHX6CLk3oVsnK8IdfrudwfOzpnQYRX9GPVhDMgzuw30+ueRL
KwMsNGOW6vTiu+h5WwJOQ1pqH9IiyJjyTMNZbYNxeGbRvR2T+x6yGX9R+NMmsfES
xnXdWNY0nLcGJ3KzgEklUw5jakScJtzoV4FXYKKTlB5J/4eYJ/PBsiqhFxSE2nLn
a0fiJb7Cr9lkEJdaPlw6Cd8akm8pV0MN9gFOtp1E93ma22vRzjnbQbEP4MFQ5Fei
vnxA8UQqRN0MFTXo57gBmkwWhJ1M7+5+miV0BsE1UT4vGGRXS+CgkEo3hrM+Liav
oHJUaQr+6I9N3UwuCVWaSlNbKmZZTxk5HKQIrxkPc6MvCHgqWU5Wk4Ax/PqifkOy
ZOVGTwzQOCK4gkVS6QZRm4WwYbLMmjpFQDyfoJLJTBk=
`protect END_PROTECTED
