`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMUppw76ZiMot2/jj7M3W+DxFj7LsYmecVcFqma3fgG+
zh6CSpExUDfDeTeArEyN1JMg+jwxwnEi77J3OPX7pkRZYRw/aDWUa8qjNd//3zzz
U5oIm5dJK2SrejgVgFDerTPEbGa4SuvIh/1hw90s9WJ8Jb3WT1bT0A5dgWSBoldS
3o3YKpLZ5nuuD3SPFnI+NC3pr0moyeqgLkA4KDIFdxqWclmIqR9u2Y7zLIG+8ZU9
KwIrBc3Kp4C1NIbUfxjfz7slzLxNTS93rUFOQb5DNCnhZ5qZLIbnE2YrjNH22VES
Z1kRvq7wWKAfktcyT4XhWWWyM3g/Yug6CWyU7tcQTg30sTlAzCdgRp4OqDZ4p2oQ
lQHZFTTS7UqjKffMJaNwvUwvn3A4BYmR1i+BhZNBBdRpCy8U5ms9Lsv5tIsUGa3J
3PPXeby+3pGP8K8Du/AjKZbAKziJwBz2Wwrwrw4yVlLZS3M/UBGDXWRAvpPPU30L
NZz4Il0hMHOdVbtupLNUlGqmCF6dnRi4AoEx8B2u5plUrSahPuJYoCS48zOfaBwM
`protect END_PROTECTED
