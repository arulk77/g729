`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAU40RWGVYtum6KF8mnhiI2sHOeiwSI/6hDqJ5mb5Di/i
ob672eBG7dXL7yuzI9agx0JtIBAOnQPotS52mL+cg0U7WhjN44WYsb/vC0O2ItzN
AZGbY+1vtRgweelzYHsD8V7k1QQlppM5j+JYqSr9U43LV7BAO/ACCJjyhtwoUkfy
aa6gYyh0+AoCuUkTpcdlRwPAmLmQ147FUHaZk2znOFCBlB8EAgdwfUekyeIQakFc
l7YTHJ0kLuFTqbkdJTMZHhV1dfOmzyunGF/TBClB4wV+7yiiD/iMifW1+1ceuebo
hzJSiK0QM+yKjmHyXLnfU83zWHPU5vgOPK0d+3WMqjM6jalQvhLqLv+MYNV0MuyX
PD/nrg2h8KQ592uzMOl3ocMWEPMdTOYJSy/Yh5gFklUx1j2Z7qSaJ4JR/sAmElEQ
ot9FV4/HLHJKZ0pEgmVQ0tq20XXR34QnIi5it0pvDq/v7vVqUiECcaUnzoe77R+3
YmPq7KkeCbAuBAvkDDKJG24b4KEIBVaU7pMmA15KoxRWPDvlcFrzbga35ObyIe/2
vMYK9tEADsEEGz84GHsCiIljzjxikl/Hj+EGHF/jxOSaCFED+rFzI4AitQwbwSLc
r6MsNgqsX7xpOBpce82CgvDDgBhl+tG0POSI+kR40bx1rTBPaFDT2N9deLB5lpaM
WB9FHA3vlqyGQEWhJsvPs9ZbxPxVhMVSV6g3Ec3R2xOuLKgGBRwnbZbqYnpN6uz9
gwOl8nld8maIW6K1PgiYBk9SNQ5Tawz4RWDer3s1YkjuupwPpXMWfZDRRwUKmIP1
vJU0PlylWhsDImirygKOWBzve8vlumxAMYoWukQZC/o9vS229olvSEvGLvdYnVoZ
pMOOvj9P8y9DZBNQ1rXQ7WwonKmhM2u6XQw8Ko/ma57TWQpF07fZ8Q4XebSY/tHo
2bnQA3NsEoNpiUM/eXG/ucSx39Du6mH/KKUFYt+FLnRVaxkAZIATrfAynvTlKjnL
6f/UcyXwPSYsMKZdAr2R/HzMt4qM8pxLikFCGGlcmb+jKKNJxdMTvnRuY4/IDd2Z
9O1l+v818qERFIoiTZjrIgnh/nGSZyjgGAY+9GM+TG5w6/+wy6T8rXrgjW1amMff
oQJ1EcPfVLi0sEbdv24twybvCVuiEyv2hNVCIPuOSAn2W7wpZC56PQFAPgOYuUBY
rQUz+t2vxJhkJH9g03IeNDklLD6WnevBq66htc52yKZbC2CpfqFAhwcNWeNVQwUX
XDQDRdf7DYwtQth6cwYq+ANwDL8wm2cdQTG0lB7M7AJsLrGe3oT6mEQrucWLoRmv
8jR/Vv8JAQ8CWsFD0uJSIrObTdV7q9B0SWzQVvwUMD8Nmui7xzFjaGboAFUgk3++
q4ZhtA3yI3+YzOYSbknKVr7VwQGf5+EOUJ4iL20JOhueyhVzRjqIL84yVD4uVSdN
H+QwYDU54Wdc707GrpygvwXCs9ntgIi/FoEG2mq2R2f0Zwrdyol3r+XY6CPrGID7
/vijnwW1/4apALJtDv8jAekXcQymuReMnEIPTrN/GVIuRM/lPzBscOEAowl9QWkv
mJZ6J9XlqSL0Bqb+guOwiys3ykjRd4QUcBOV9VcUv+WAb/Md3rHIasp1GSX5fleY
bm2iGBzjm0nMSbvtr1u5ZOoLxHVYkzZys44Tjbrw033CTEdKR0siztdQmCCJT6H7
0Pm/P5HrZQxalgfodnldCqDCWy8XUlnPbZ3JiVGv82cLa/9JUvpHp2dMQMRv4U2Q
+luQVFu3O+C3O/iGPyXD1T6eqOUE8wrXpUFEb9Ahd1m4KPNti2Fkx7by2MunFtvb
I2iMOj9AhDRP49gu7RbEkvZf8cSHhdUnPqcFjPWyBnArJ8EM72iViRygdOFsrzA3
lP3kzm5wfsX8fx1FPFFycp1KHwxzq6nMLigNjaNZwtL5G5tsmu6W2I282fSOqg3T
jZQh2fFD7t4l4EeDpIXnJV/rDKuYf68Z4Tq7ebwMwZUWDOEUmIaMa3whyzoQ2S8V
kUDlmsWqfTjl29AhvTXtTaDwHGydyyoJxIlefEAFD0ugHgxFv96GiBQAt/qiyPIW
9QPuXSomnGmfUtPKZFucZmYZdfA0CkNHNjWoQ/xM4YCMI2sI6f3taAqZY4HzuSBI
IMbPHutIw2W8mGSmeN2hMfdkK2BDRvgjmoQIzGtMC2BY89TGbaNBYoLiQtQNbYzt
2GLvYW+OojHW3FO5is9DUCDg4B9VwojSNv4ZIe0audhv9hjMzGcOO31cz4gDjiZp
fjBGUClqXw4/r2bT/COMBK7wX368HvalSNwE7xKDYG2mnBPg98yJ9ihsaHPjACX4
+V+OhxwACytDi4HTusOjPv0Gn7PanflNHLqPSkl5etd2cxoEzfrt7+ho3usxxpKQ
l4L97y3WLyEtQz+KhH9p1+fxiM6jal5uQVcrnh2XTcMSpmg85EOIHpjBkB+cxrqy
JJNohccgyjqep/Lcn0C6ZOYILwDRDcAp9SzXxJ8vjWHXXgUnqADRK1VK9MOlt7oe
zzfR3pIcXhBC/V4Ozv2EMokPLbOZTXhHC3TlrGTvbLIp0ySs7SfBC3Zz9qZm9tl6
uyrBWinnPCG+zs5qt4Ml4mGoKd2rgqcQQnCsluMh24mK1bUp6q1osiX0xMVPY3y7
8ogBlZ1fmOXMdMDXqEmxVC1hGouqfpVNbvdYDEDYZvhdFTXbbq0hU2eRlIS3ywtp
yKYLV0aPqggZjvrGxSJVBu8/ub5cT6INz2hBVsJhYU0sfoJ/vpjnXURDRE9LYJt/
FEOGf5cNE+upLBMtya6rwb6NKygue8lqdstTU/3qQF0HIAW1UnLylGEQk8TjWlc1
OtzxwYkxnYbcJfzXaeCYLmnW4EW3dNW40aE6UMQ1ZHR+PPvHM4sVOBY9b/d1RntQ
l0rE4A98DOSX1yuAEEFo7E7UYrmyEsso8kEu6hNNP3SWyV95QnnOPDN3KP5mmnjW
WJyLr8g6Fa5IvKHn9Gl1Sub1QHFJ2kDLtl5h8mfduFkqBzAGI4fmEBLmE+JLlb25
hORYqKfgFbuoVohuBatuZC3tRb+3tRaYsS7Zt/uxYSCvj6jmQ7WPU27K3dN7euTk
ErKmQD6q/Pa0/HjDkViVFzEGFnkdMdpjePwajlHvUjzeSAHNstvb8C/4cmYvEhUc
AhscAj7JIkIOH6uqA/4vSjTeJ/SB9Nkyhp8y9nW/6V5ujTrWMofCqHFMzWHZmTdb
Py1Pz/IMxzTh9+/42bBUTNVv7OFD5bQqDLR/B9Bn5hzK4PJs65RTp1Rmw3Dns9U7
paDy1kDgm+cS8XSdlkAXN398ou53JkmLGNdy3Fwx8xH/hVZjMDzTKEZsK8yqz8wO
XmYHgsa+acNvZi6/AO3j3UVqfohBDYib6E3g7J2eCYhnWSoMEKTsMyhuIarP2L7+
ywBqwmOfogNvDCbervIB4M48RPqcYoEDk1WpnhZv26R0ou9XhMKXGObgQWBp7fWP
7zLv2a3N1QtEjtz9sj1P1J8JSUcETydc/csgFeQuvc8kU+kqAi7Mu6z6gtcOA6W4
lpGmMm6E0RmFuDV5msaQGL297CP/DA2JPvl65TFL9jLZuBt7UrvgyJYwAqh+SuBo
Mg6UNZALRGhkl4oWjkbwvY9xz3Xoxdc5NWU0SfrTPI8ReXG/QzwaDlsGtnymP8xC
O0QCsYJj6jIUBG6m0x7Kf0840a+KQzHEbNtjzMvgumTCKI+YMosoXwkDnb1VU5t4
pimVn7J94gZgPxZq9SxaIXZbBjozZL/PLhWnnQxw4ICjsqoF19YzK5NUWV6ocs+9
ixQoPz/CkeTN4jtxpA5JLKMj5AmqcR7DnYHfO4meMtNyIrQdzFQwHE+Vva+KVKTC
WqlS5sSl0QXM9/dCY23krRejFXBBrKXagkPcJ3MQrryNX6xpH++1pQg5um0gG+n8
FpjZ2I026NoNMWSnhNZgnvUQsSzJVuwxpSDInn6UWPflE5f9JcZaiGyw8G+bTqRT
SlU2W8GHNnz6IsPQCZvXOHNOCq4wNZEgmEuzeHGBPRPoSQXuWhe5lwVV3z1rEmWd
ceHzdDg8skorQapUDqmoBnS2use0F7KhGP2nz11QdJLuMeXBfXZ4lskp2EGJZoek
WRmi/1lxceCRRUJQnsqspvEOwSjJ0NijhSGuFG0p7bSa/eGCjoXuSbqMx6FcBovg
7hejk70ll6dqsdXsID6QRKxequetOHacs8w+xttkQ/KiAKR6EhoJ5SRdG0g5v55Z
XeDtQmFzfzn3izAX8r26jlSkUnOVMEp/f2p4NljJdFUu2MhpRpV8Ni05o3HxdJaP
7b3wKa5rK77l7GHUpxP9s+Qw59duWo4YElS1rcoiRVSswACn0HkgAxa9Jd3eRjKy
+t4fQBBJMqXoW5mcATVvLFBG4bFABqYSH1vMaFo9ojYOmAaZMaZodfbhJD6SIFQe
bKMBKfy81DkV7WMx56M0ogmyUNHDV5lIv5SlGcedU3Hq84gw6CSF940scV8+icJ+
0dDY1hQ1qcYVKlp3M6qkYVmNB0tp8+pBxBl7P4o+abIZXNesOE7aBq9Iq7KTjOhv
hodmHQssB719ZIqEYV0mynwHXhZOzJB3CXe6nlRwiGfPcCM8CJsg3wnlUbOOsOmw
43VGhtPbdqv6JInv7dutfxbYXzSIOgNOsMtw2nyQMCeWYAVAI7jaE1iFz6SAGzwZ
DL3s75jVg2zxreClOxNLE1Zlv3HrBce+pbb5U+39GfUD6rJ8J6jusE3bmFvcrpME
PIMxOajQoz2DoKgDvDywFQtvZeYkH2fD1JjrGJMYUbC+5cqGkVc2JO8d8XkSSgdh
esxEQkf/VTLc+gOCcNaf+orRiAHiwnRiEiiwSE/MT/tPBxzPNSwvXoKwKuoQHjRd
3l4WxLzAgEdf8wGMYhvCSgnwjzY4xgTZNUarUydHY6Y7e9tJeoIvvdLfE3P+F4/S
fgE61lH85zHUDyu2+yOvIfmqFN7bg5/coIwydEw2yTdTdRUFW2zdMjoN90jWJ1wd
xC8+J9CI9e2hV56lMDhuz95lxZeIApC3FSwPIgnCJ+CmNRz2aAvUpMvPxljJ/Zq3
oZ0DH/gpMHrRbJq9+jtbAO+dwUWqVcpn2ZdSR3OZhThC4tqkFxNzetJt8KL8ItCT
AhmzP4RLZh4RwnG5dP2B0PsrZfQQN6glIcmpoVm7PzFhhMKXF+BJV8DHSEGk/xwm
zF3caoTvvwFmm3ZlQ/MKRggDD/W+YJgX/pycOqzS3hUdaY6apaafLGYHvvOhfBy1
KgQCdfNMeY6Z07tU4swvqLL59dwV+ReyBqN4G1amomwrHBJ/lSW+pkmgyGulnISG
2NhgXWZe1Ama7ugayXQzE1dv56V3W2irufXCya5f7UXPsp9AbaP2UvpZ2UGp+kT8
3NJbB/251fHnDwDG+w5yEOnUyPd0pUYOuzAb4qGraU/VNtSXeEZqLuMIpcAcVwul
Z5cNLpm+0+bVI1WtHT+9bCYjFP04LRa0PGt4YtKXXtKK1O07syilPCFmih6VN1l3
bDDMVCLYrwab1RsXE+vsgcOYdBxhxMN8ZplziZgvUmJu6RSiKHgluJbmKD+MloMI
OXYlCk/pr0ktnUEXT2W7LIZwjpHqSggHdzAkieJ9Gd8KgKv/JkRoS7AytZtTRjR2
RYXQKYoef8EnniVS/q/jHqNk40cZvHxv4Pfm7vHIt5p3EwZ77Qf8ZAp4ogw3KhMN
p3GBZdpoB3qlN8PrhJDwq7ar0P6oLQP7h6tIcMsQ0RcPER26iwFF72d/13Pl+euf
miu0ElXLyGP0DE/Pojmh+knlEklJTnOo8DjgTnUxRKisS6864o24OVatAgNKDL5Q
1Gpn8ne5Nc5RNz9GgHVzhNObx8roBFKWH+wfO0SSE7L7J1hWnfbX4nvKprsJoxXl
LiLT+lk+t33dZuiCmckV4AcYULTeVtnZ5ukEzL4J2buCY+LppKu4j51eqq/ezWRN
pldlyH7HZkJHX+IhMygBO1eYpwh7hL/OnNLfa+ACmRrOZHTn4RL1op8m/x8LKWda
ob1uK/ZNNKrrcEXm8nUsnDSyzbq8Bn23G5xHLWk4ZQsj6lU/JNn0WPJ/Bbp4tBe8
pgVOka7EtHv+eCmJrNSHMNUbPT0SBEPEC8qqpKU791OdoXOZX20e72sbfvQDYPZt
I7F/dd7PazFRIQTxzIyJirX1M+C6GNvs6gLiBUubouG3qx9sfCESGcz20B7ESa5D
XozlSdh0fiWGMmp5clZwb6D5gaYWOCPmI3zdtpaqq9rmvlv+tdEWq1DpPsYbc8wY
7u4cohzsTSiMDV61PUXmtu3udatl2jmoVG4H60MuGZVvK00gf/muyNppAWn4pGSe
GtyqGrTweyfdt7FmqVoCw+u/36pD5n3igax3D5sssFAowGFbVv/SXX139sXuFlaq
EscDevJks/VUY3x4UNhlfMSKGhcw+btY6GIuFIO2BHEQmDt+aGRmerICtXlytgOl
ly2YLmUeAAz9yFI1Rw+sV8KGrYeXgzUU5JvZlcpxA9MD/M0IAm+msjm8gnDuGUOK
Q2Hhy2NVIk/Iru09fr58Q7mE4+umo0Fw3TIc0rPVwZ814zQSdrgQiGEpNQJ6N3Ob
tIvP17ONU563z/zqFaM0muP6LFpT7FiBwB/W/v82fE7dIqyVp2kfpeLa4bJt/vTI
qwLpcZ9eM5AeuOT2df8VKQPIbaAr9Ax0ELROt30oOiyl2yySQe4WvnRLKVP7RbVD
8GrwLnJtFqQG/itQCk+BWQ==
`protect END_PROTECTED
