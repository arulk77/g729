`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNZ1FulPzFWlGkMZmIAO3a/UC3xE5YyBqxgH9g3Z0UVQ
XsXwoLGtOw6RyeIcaLa97LaGugHWlduPlwACyaghJL2oKSZ23ct/9HlOXzt4Kxbi
QRWJaygSf88EdBwJY+cqUxgUtsKmzOs8jgldsy2LMMMUlwYGUUXj41vMLsXLBsq9
+DQLpRZ3iUwMwp8VgGrCG1lFuVoXRvWtkaLv4aL5gGugV2zEdw71B3wJ7utEdyL2
`protect END_PROTECTED
