`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
s/aNTlGuWifuLJiJgnUdMdD707q5qX9ouFHtBGK4JcCbDAJaAz04boxfizkEcvJq
NhVTwRd6+4/kX3rT9tcuQNMlTupbIo9eVP0ut3gxaixXBhNHOsnNbOLhB39CYJ7I
EZ5L3mEyPJLAqOHTYmPzLROEC3T1bzDk+gZShxjI0VL0jPN92Tnx2VN/xuL082Pi
O089gbrRAwcMOlv++S3i+pvLF4Cqg90rHOt5Rk5Q3e0=
`protect END_PROTECTED
