`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveArUmwjPSQF1UIOMpUr3M6f2796ddI8LMxjk1hM6I+aP
XVTWMXqBCNLrYgb+XliYDXfX4pUKiW1rQUr7QgJk9NjUN+qcdllK0fcYuuflZLLX
vn1SLpisVi6vdYB5OHExXlW+KPjsDGTlVY3CzBjXq0me1CFnLFdYAzoXxnhVRdgU
NTfVclkBeapuZqm1FrN9u7baZgyWgWeA8GluROll/SWDflxpc/U867MXLHwmHGEB
/G7F4VlbPRRylAIa9V2+i88ral3cjJJwf+lh1R1PlcCA+1y0K2rWaSSacHEHOB+J
soQB7DiIwW0zs+D7xXl53NkwA0SN1FX3hYX82jY6/OWcbjbCZZqJ2dDtqtBBo7f2
`protect END_PROTECTED
