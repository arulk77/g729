`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDqBmNKGgy8pJ+bWdSWRqSER8pNfJZ2Q1FutD0MN9T2b
3TDw6SpJUUvjQZcxwqCj07cpwFvq2/VPZaFmUORI2pCGzrhWL8fpsuQbXNmlroyg
6yQYlGeMdYqe7DFGqsuGXwPwUrF9StvRR/CisoORFVH+YSLW/OAAkPxYBWaO9O/h
iSgpjyBLllgXuLFhuWOXqjc+pO0a18CoaYEirZlgEQRsUt4YdjWp5p9kbiCtirVp
90c2F5prrYxGzuNVHZDVVgggv7m/cr/aXkyOqcTs+DLuilxWuutzK4xVR1NKDPQQ
YzttEBdW6LghrssZNLEC6PzhXZgCBExZHU0MFDfPEqCJtJ7OnlOu9yjYgSCHkI2k
26uALq6yb/J/vKznmiTjeN6Qnf06IuCtZFWUcZNdUIq9ZglDI2U+VXRARXN9XroB
kXbojxc3sZd9LNns7eXCqnKezHNkEJBCH00sRNp2PGkcHX5aehAEzhaquvKXef8e
hfFtFyGHvxDx5IZEY+xoRg8Br/OafZrolmyvWD9/gTDEbty2VDMS104MPx1riML8
7nCQxDDbl8PZA0EvUWrrt0RgsozzhwF0BM2yg7SQfzQroWYDI0yhRmFe/nxn4Igm
IWxUChFRkC18YnGCJKr8AIBbSeRqU0TmnyIn2sg5nBKgZs56vKDbrfT0Plta9Puc
`protect END_PROTECTED
