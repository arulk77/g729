`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
wxa9oOG34FqZzPEw5tB7iI3i3i6wirF3Xt8nhdx2lITCcvQTNekHnaMy3XAEl2LX
MW1tZHBeIoQVo1FnWT8Hu2AxRHcaRe1X/KjuvJcmwCZ0N9e3oZE2JjviE8yBsUpG
OYP8NQpQvS2mDNguQWW2BwjMeN9RNRSpl+XMgo/h+Xa0AykWOaqyivDjsiDmI624
30rboP2LpGCKU3uLQeo9TVmHpl/FAHLwHXGMTc3efj/aZv2ADmVegsRYBeyH5E3G
xDMxCF/0ppK7egLv2V9tU7uKjRGpY63BRW/fnElP86V8C79EE6iFV9qDdlxM7paH
2peCq2YVpr0QTt5aUFGlnJypjMXmQcstreT/4FvtTz//RoslDNwIXlxYjq59+QaW
4ewwLZrjjO3gunDJGyA4ega8AF1nZrK0iJLmRcNYQI0=
`protect END_PROTECTED
