`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
HwN6LxG6KyNm0WqMHnHgil3NExPixhcQurAHx8zPdmkz9t62R5XcnV5bWZ3fxrG8
bJg0nxUiJFNfKKzVyC8yzsrsNq5JvhI4Vz4FfM5ogq2kDa2kDr6dZqis+l2NC6zs
7NgLJb0EhNSiUVNBLcv3qvtbqhVswYDhqMZoLd7OOpw7ZeJPgyCKFsNy37M+iEua
URf5zlDMs0kqtO8jK3srIgh4W0IWACt8gObY8ksSdciD4E/zvhrkh04bvD+paEJX
JZPTzH5RMnOw64dXkPfiqI59K0V2kQoIH+6+bH0ys9ncnRddruaBsk6RfG1uYu03
zZvzZBrstnAzph/KLuYJ4QUDpU/yeVdITlOHin8jPDE=
`protect END_PROTECTED
