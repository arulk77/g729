`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43c3UvaLEf4lxPuB0lPvNxRnRP9vA0+FXkcSyUKNkdbc
ilPEQ3JmWquXwfWhEhIpUIc6pocRUsaH9dm0ayGkm8mAkjJHW/1ISAsrtLQPdppi
i2f6WwITXU9Jyqvg3RIDTZUG1BnXGxFSK+FSXLWS81IGCnaTUlOL8yrVwjiAeYtp
gpuvWRYl2HEiNgFia25p14baYV/ElBkV81IGdvXh2wh7UxUQ0BlTL3cdDmcv7ZXj
eTurMdQTNNwhQ8joHT71f8y0GYj1Wl9qbG1uF0mVCFWFKzBgbI7N5w9wZFSOiSJi
8VmlgqywWrgER4fO5k6PwBC5hZqEZtbteZq/smMz/nYCQSi5sS7LyDJ3DqBweoLG
PYMIVNZMaWMsrhMp5aBWkWiuNsCfwGtnshjhQpBqrmwameAmdPhId0QZiLYpu8Av
HlNIdV298kWJUSEb7YM+tfJYU6QGIaclLtgQUjWTRdpN0EENtI2vGDbmmKuZ0kkb
`protect END_PROTECTED
