`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMY9nAovyctgr9oa4n162z2hy1qegDuDNMfy6Labp0KF
TKoy7jl7Bc662qS/bBlugWdZzLtOaLVY1m/39Wo0odyMJWYpNo8rvRMRBAAhBOsl
q2nTqeC7hDXptmxrX2MfiOQ9piOxye8cvqO4Yl2wIDHoI3hV8UQv398/xt6jO/Gg
4k28uXJsLYhuw2Yx/iXp194vBI/6H8HELvbahCd8BMag7TI4xdJkytx1xxfyXkz/
OkVPESZ5fbpijXKmxYHBkmRrmHIpmkRJ3W5NTc6wyQugzlsMLLJtejGrktOoNj+1
Avttqu/kkNlv8FIFpE6iV9eqByyNXXSLgQ3J6KQANttBeLeIwo1vVwqx2jnhDkYs
pcGTGhAPM8KT4Fy7qAQSclafB7SYdLLpMEOWp+YelMxi/HF1aV0kDEhQMNgh+l7u
s6FoPvYitQ+N4tI4XEU8xGvzkN9YSasGdMugjVHHdHeouCFXtyaLV3UaVmb/WKAV
ZcLsoW/eT72wklG//MsuRejgvCkqanUNLbSEATUIu4CZFk/CLy3geneSh5KW1hgu
Mb9qQKx3QN455+45P+Yux2Gm1lDRYqXOiJ3QEtKGT3RYG1sczeypBesOD2f3fe3p
oCz1YkFhxCZnVtOi3kiYssKz+K2jaH4gNGVKMhw6gRPfrVWd0KOjyINANP9jdWlk
Np4s1qG51nRIfpTwmRoNQn4zxRKHv4HNDfqPzS8KaowB98qV1MuwxtKmm+1gXdwJ
iMieZ+bdgNa7AfA8k2bz4egtWS81x+E23M7hdnWxe+KQ/ZwObLhBeeJ6cUBd85wm
AnIFR9ycEl50xjXxOXDBKvDb5+IvCP9JkkeTnZdCxq5ZK+N5aCKn1rwSFL1TY2+3
PwEUUBjx3r0SsTx0B+GSECBr6Ay5MAEZHX9VIs3A2EKE+ZXDdu7CVXfz8cRiHHqv
IP5QzzEzeGJeRSgRpIzBoBlxRduFLRIC362o9dq87/pBQUM61V9H+ZIEeWrX0MU2
gmYgcdXnCLH8PY6m24G/dDQURnjHj1Wicf9lyHc9uiH3/vvq/XxbZ2wt4tOQIfdJ
hEcyYyR1/1JblQuqK6lDRu2OwxupQRlQNH+xEwBCEvsw8ZstsWE14PZMoZoD6/ej
NyYw4xsw4X9HIsjFh4FG+2XXV50PbdSsrGk+fguLM+kUeJPzh2LDOnPsyTONMAQP
3k4MRM30WXh0Q6xL2JA60zwOrKDPA2F24sYdwO6aeDqWaP2ho8denVlERvWF7dBZ
a4lXTOtO8KeG501OduMdCxiiRhMQbcWf6lppVnJiGP0PhZkXFr7z//FVC8jiFv4X
rwgfOIG/LRAm4CDyMh9jO0Is1cTLqwVqJtz4vLbW2fGgQIwQqulabILaasGNqOM5
rQgemSVAMBzH9qxWhhVDmSOjOfQRgVkD8tJDd1v5dkz8WEJZBk6NeQVeURDL//65
YTuyx2F6Te0vK7Sbt5NxWJcH7rqEcbaXQJAEazXNRi7YMK7zLcCwpkyIGF5gdoAf
aqPUuhwhosnQQAnYj8uRuEfRA4nrEecsnHUoN5XZ2THC8M+d10ALyYEI+yNjVI75
d1BxgW/8EDUWjyGGfgZCnHHvkB9DhNe9s4tz4lz3hhtomeaOYz68O456mKSgCmdW
nnjKTGJ3ZOFh24WYIhtV04e0THyezgK79CBHvzaIMJ9zPfeeRSL3VEPINcYG50Ra
8WqxvuyLWSeRcKYt170jHXHMA7AmTNMBuyWEAcUoYCjQvAVKbnvpccJw6WbuU9lZ
ZjO4s/dpVPPgaXzgmQWa+C5tRKVOYcjeITB5aMU3ZXwrJUzzlE+Vl8HAvyFRIPzP
eCVb+JtrYkcOR8FAwAMhL9djR4iBGynF5DuH0R58svAkbulsGg2qkiPVzUuXmt4j
F81IuctKZ46g3euofm61W2QNNa/fe2caPwaBJDCWv+69ys3YhZ2Ytz+8iZLkTpAt
mwrkuasp4VN2tJHt3IEbr67JY+NXf+anGgKf7aXzImJrivIdl6MdF8PrbVWwd4X2
UhNs+GRXAndbSXsLDbX39wdM4YqVFRa5Hbr6qVpzD24VO2pTEHP7FNySskpXD4lS
faK7JENT7sdSzqCAcYRnsZfWJTnNsynF80D4PZhYVCgvtyE+UMts/qaalyET/+DY
N3yzTPLOadwBa3Jmzym7lSi/9GXbdNFCIhV7zI/0BLKzwrllY4I9lf+mw6xbfQbL
/9tX+AFtr7rIL9twApzJRLcCNGiVjLGgqU7PS4S7j7K5Q1NgieZrbfQ6wvmuj1xI
HY9YwqZQJJBPvzijBb3TTX2M1iPq2fBPq5S9f9lFHd6pWF4EDe1ajyK94RmXWr7N
ReyLgQsfZudwT9JuqiLxNBNXKtkMdXZmG2kxuJo/fVtyE5RtrKP8Buppq9dWcnsl
VmPIjWss9Wraitzp4sQvw7kXT0YB60q3xcqUmQ59WbwFNjchyRyjov/2PoUHH2/9
d2c3C/7TVSRjIQaHMoHM609VIz02OOolHElgk2o4+NrWAxQckStgpGwJVm2zZMax
g73cKvzlBqQqeXe6vbduOAjzYdXbTdGukjpwlYVRnlsy5RhpepoeuxRQVkpVwpzi
0XSNdrEzuTVjFBMcQERt5l3L21gfuZ9GZmr/iRgKCoecdTCx9fQ0nifp1dtDaGKl
jxifdbYGgj4U8CPRiZN3dstACtzlfazHDIHacVYd5T1CBUobmAoqreYwGuISh/QI
+9ffcSSSA/t+eg8Yf+rf7wTHEcWAujwtSsf58UmccpTzj2iiiiEuUbcFWfEqcVXX
mHusY4ytryDR1Dy0DVf5HemTKJkFqS2k+j4aLlPuHg/+vAhtho/WMldzUtmXFZqD
SAx7OvxJGcELvEEg8VK7NwUf44ahxmH2XMSw+rQMDIC6VeaCYvP97E2D3QKrBHVo
WDGwIcxEWqhgdsNG6I8iarhPKcQx5OCwnekWfM7AIN4OtnBfBEQpK6G2i6CPBnCC
I18nDE/t+9ndTGcch46VczH1lfd9iLJ/atK6ma6O/vQMNj/vq1t6EUmXB15Dinzs
JDfewNIHDklChHlIeCjD3BH52oiIFY8wfKpwtUporjZ9Y0rlaWTho2WJSRMk6/tz
3qQf708AUGDIMsSo3VZ73SA7UQjBZqaE6w2FYBNfDWLfqOC6NRyw4GQOggBJrPDY
0+K0X1oJ3E93xfrICezV8kbQpWLYxqoDXKg8H5ajnhr4EpWQB8XQ2hji6VLXq8+X
u602k0zBsroDQTmzKfVFoAVVC9zXXCDeG9kXZZXA35DMfehapNvE6TqnzrKhwYtd
jWWeSxjoJwttytb/nmulU/xAKDJgB5AHT22iyBe6g3XRAfljrLBl7T+akOOy2qXb
aH1C6/o2UcWHzCuf8pbVFpEtS0PrPJnRtnoGlAYnS6emyTI0eQGMks1XcTUKKKQ4
Y3tFBMwh06v0wnnhBo+hxF7zgGeOP5vpZN3z8MmT3xbYTdFlvAbTEGY6LNmO+ues
uIb4GSXb9eOwzSz5KWTKdF8FrH2Cvl1w27vIApYtByAwe/OisyORNVqFmlIZpKNz
/V9D91B4R8bK0py/mYgJ7cjJQsOCcCEVZhjN8627K9CXMsab5fpndyZ8lwjmGl2T
69mZezkezuZt8ZDYPKbRPBAn8tWA+hRKvCT4pnTKERRV2KFQJlpeUz64bdv6r/0H
i1tvhlyw+3JVU5X6oFYMB1wYg8o/FpgnowDNcxJNRwRNhIWypHAXK7TGX7tJeHa+
9UzixN0g2vGzjyqRYK4woBnb605N7xE0rbiyMgehsXOTkBhFRSGMmIYGGLvcHuhm
rA0yFLw7RTomnTD7P8OkJwetdSx8GwqS8ZKCaA726EDi+ouSoSYeNbu+NO9+Mmz0
+wFl184KUpp+4tQcmV37EcIOaxE1iE4HbWrhmWgVqPR7knOPEsizT6mFzJ/xcWBg
7Y2Y5O3LlLTX0tX60foVEnsWuLtnpVgng9O0Uo50JgZXoP50N+QfoC3O8XuIdN2A
7I+9/yMpBC/6h+SHlFDqjYXvxTcB4LEhuSJi3eD6wASZUvYb7uRPpd4y9ARiU9A9
jXDTXNQr2dq2047FlxxyzYNiAzu9VDZvgveZgpEVoQw0+vWHnIoXtI+kMuarBsMl
/8Z1G6ULTmydLDykzznJpdDxee4tMU2v06mgRZwEZDIVPNwqPHCFVldKl4NfzeRR
CCjR7ljc/MXk5KaiyYBZiFEd39v0mg997x7uovuU6KtIB9Bk/cY82ldxV6OYwy1N
HERYEyDsmI9EUuTwCXJRokWXorO2dVi+jaPIVqHolQi9kPtW8yjXPpNADBMomcR0
E9sfRda5cObIThrzuoxWqqabBaUIvKWYYwjj5PD/S7tWJq8odslpAicGMzkHoUJ/
b283ZI0cs3+VSIkgEV8wZ8LYvc6dLc/829WV/AKnWMuljWk8MyGipoao7xL6alkS
lDxayavWzWPk6zLW0IX6DmAjXXgUw4Ty12RKFutlr2HqQxTb1h57bbr3SYfyY7Wa
af8+vdNuGkxGZW+l2F8hLvrj17UCBqsVVDyd+6jtS887NzakJE82iiLZRClGMrzP
o3G1LI1w47Eq7SZSmupaYuBnqdyI3+iwDkrNE3FWqoGo1I92IGql57ATMLAbL0pK
Y3xS+MWzalt0b3knL0qbYZFivjvlOCDlfL0ojkmwgd9oQT6ayZtz+Rly75KOcvfC
HSyl4iaGFHMDNGu8lSK9QOPGqlm0vgrAoRnDASFqsvbbq46XBDaDTls3reKVhZ4p
eWs4kzT3y6lwem9PlNesX9dhuEmGiQeqytwGRsEe8qoDB/ZmjJQChlWbZ5BYMwbY
6Tb40h13rpsEYhSh/CSufWWM2g/C4pmDs5hz3EroeCrqSJUJv2R/2XNQRhiknNvv
Kq9sdbS3LaDnbnpb9Coea0DxRZ1r3xJCfPTbulAogEm5AcouBl7HwaaHxWRJXFlS
J8mUyu1x937/lQQw20AellifFXkyKTqagGFT9//JycYg8ViMBMbyckBIfQHH1IoN
mbwM5CUcg08NqIw6oaHsd0GKD/MAK2bgWhN+u6Cj0XrIWLD88Z6rxBI0f/t3pVEE
KAKuYFVmC97W9cIXlwGLbE4Lc7mLk4JnhuFZq1PlonSX+yiMD3f8HeD2dAH1Bcug
NWhVLpT7NDUDSw+16rWb4S10kXdLJlXAKrpWxC1wX0PBHd1icsuVD0tQ9oNjf0hM
3P+B7Wvf4fYJ689Xmt5yVj8/KcB1pOLDP8BlRe7wprnYFgQ619/bZVFiwJPXIJ0s
P0TMNERTjh9wVaoyGRez4hl70C+Zv6DDoWnhW8Ct59hveeCYDM97k48rgoSOnmVl
e+rX25ObsHBe0/vaYEZs02Z1cChcEiYagCzjdrZ37jbyFGnDovzC9onWLOT/Fwgk
xv8/mQBNja2JYcSYbzYP08rkn9h7xwC0M//D7TlWih5SBIszS9NR/fDCe5UhmGNy
PTn5RxM/RpXOrQtOZbiqBvUCq6s77wz8ysXloyzVE1LEST8YcNshuJj5vWwK2PvR
g0ZAZfU5yG/DF9GRKhyKcNGC9eK9tTmRiF9MRTXxTQ9dLLojRXIVNg23O5qzklEx
y70aq1VMgWrLtaHwowM9myOwS8WFmqANc4ovs6xXzv22yCkl65bm8vp7GYltgJsy
WVTsaMTByOoKE+vu62uThUU0y1KFndLgp9AC5uuTaFoT3dCnpuF3bvPjV5vnoHXk
sVnE6BRiXerRxAe1dEeLdMBfnIMqOFRQlPdyUAM5EFmGdKEaxNu9YXTWmvch8FPm
5YE47x71yzvC1RqjFG/66U4sfEyaBdSQh9BG1ANj7DY4QpDpBRmVoiYp78/KvmM1
jkGtbTALeppwuDNm1J5VWLcOLUOx48pfGlHgIUGq8vcfnWxQhPSLRTiIIaAT6Eo+
/POz1E6sXNEFbxD29RikZEvCmGx9/EAhkt69WnxsKLN+yN4eqmW5Oa9+NnP/qsRf
d7u1eyzRH5Xdkl0drKykOVHXW4QeXbrnp7S9GB4PNi6/d1wG8K0klmcHauDgLHXa
uH3eLq/vysWUCm100JJ0Ddu0cUvwn843sd59t2XqcGB/xa8FCkVMW0Lk3NqPERYi
OE6odYJsLXGm+xKnzjc0BlfVxrq889WIwcfgsDE8hbfXfvBE3LtliG2rr88aMY3P
W186KfvF3c4njUWZz58EN67qQBVplzZ8nQ9FRwW8Q80p+XGFfuTWV0ImAOC5SQpa
iwiP3rOL177hBR+OPcmT9lDNiJL8PQl9kXF5D4GxwmCDlMgBQ/GJn1mAyPkNJeOS
/4L9g6NmUtOLaC01Gq2eOjbinP5cJtpA3YM8H5CNEuIENV53Xn5t2DIB0HjOrW1A
DYe8jXSnq6Pvgptck4FxQjOw5fa53iPZ12IVGh7PN7z4q+iS7zV/wpONlmvorCjx
atGvqz1rnFKZs4WPSHeNdHnyB/LsNwYrhpxHjTDWe28PBHsaBaNq7CHWfpupVwjo
Ej8BptQ7bSIRGvcPJVn1UaQ7GfKe5jugpn0vGhEAPNvj2fMlnmLbb4PM4C8r/kb6
jUBEy/PuJ83tOMH7m1YhPrB1sAutpnDLTMsl54z8D57tPPMAH1PkoypkXe8OxxN1
3UnUpfgS/vVmcou5P8g2X1QJaHBm36rBw4Hv7eGsaorbg0z0ozTMeVK8JcieqZ02
vcuDWBlDzam9Xx0k2GOUZPZObzQJGbopjSMFiCScVQ1y7s2efL3dxazQnreG/q48
okzpvvvnMYNOgY40T7vXdR3k1d9EroxC/MnZYrynEeoMzrCZmQuDfhNeUmEFhzG1
5CG0ZUK4r3Po4e5/bZlrKrHLosTXTgrDYiuKgiRWVsXi11PHPx/YgQk29Miy3cOa
QVdT3Ng4uJ1zP74TUbYNU2AVVO4qZERcaH9CSUJno5mSn5PilnD1lXXOvN6AlOZQ
uhnUdB5bOb5F2cdO20ZsdBiBw18ff/ThLyVjZeIQQdG1ARq9g6i22tzKT5qK1Czu
BTi38XFIQeVamjR+g5m2ufosJChpOG6CbvgyPQhM/LprLlg4P0BdxePQdXNZ4VGx
dC3rn0B8qhOdpHt2sqcTULeBf9IdZOxS8fC9vOcKuEaMUcEWr+Nv7d+sVtktd5sM
Inj4FSLYpqJHqhhRuiMd0tCK6WD0SUMmKlNyyObIGLPgETtzEDK+B0LEGc/uBK6V
HBbmHzMqvoj7/YtuZ6dtJ7fFHpfb9E7hdxw/1RKHvEKngU7yaYaofbbeQE5TiprI
bVwCHgoIA3KrbCUrOvOc5LQeRpXYZtoipxSoN/f4EHOftsj2kWWm941dej9hzYMM
bkkuexfeBDfwIOiITLAJhODtIOPueLbAHpiWCxBiEyq+mTKph3eal6HqHWkcknWc
Q4Fy2AMzNgGMs/nGoiZnzQGBj+D0yeeySiOVfRIBvbUAIvHBwbjai+gfEyFAhSHA
SJYJPqKXdeoYMeJL0QsMjQm43ErMoqatgFTGMKqkOfxSD08sOuqDOC710Z3HRfKf
xgg1hQlm6oLMvsvU7WtOfCOZnGMY57vqXOSllfo1+od3+JLiIrRlM8/riUMoT7LJ
rLGiTPgQWzEXgaCcFnX/i3+jFg9hGTrAjBh759C1OJoUnLXHMHCm+yFlOYp/cQ7E
7s34YYoLjinAbMqodKV+yKeJASvSHm4lU0Bs5+DVb4UoqZBgutUyUw17xm8+KpEj
Wg9ntavzDHSNTrQlPGwtKJLrjV0c3MlHchDsYql2pXMwMxJpXhS174IA6576UuWR
kLymhZfo6J1haIU/j9Bm6w2E//XHSIypcZK5CcEwaaYyPI48U5FJkIxXYqOCVOK8
Kk/VlIzxYl4X+oXNsE6UAdmzsvp93r76IuKaFycWndnl2PoVO3EvVjJ5+Jahy2+q
xg8s6+v3IcUl/czyOTjSy/Qh9m3Gw6+RPACDnFag1xsOsU821CgUfByf6fwgZVyh
jVB6tZbqC0MPru2t6c3d/axu6d1Bn/WD0L/DYTnXMRn2/1Re4wQE05wqY9vjQK9B
8EoEfgzGZ6jzLkfz9PMI6mjceoS0XbxgrssK1D506azpw6/g9943D7CxDlIos0lu
T6Q+2GxsKWYGwe3JgQnmbvPqPJ1N387jWKfs3siSXvAUkZf5G4tVtmRXSLjgpX0c
tM06SBc8CDJ4J+SCntkyNIIMYBaqMgsOfHz8DormO+wESAw9mqNFTTy73jcHCqVP
DHld+40J9jCwlqymuDLRDwobwmm3NifQF8duutXMj9IxURQKCL6FuPWF9+Y1z5PH
CWto95F3JaHbXfOfM2bTifY7TN4ApEqd3uKPjlExl2IRqi5cES+SVpF6MtnZmool
triveG214mdUFNS3rKkSpaL1OcpbdDBKaBbSYarTrwO6HqqeW0nKSYIBo5pvrdhW
jRa5F0/vTIG1GQKyzDlKGhlVJq6oiToiBcNWEEaVcqqOIvduiL2s1hJxr0cmqYTk
SDOsVutvYk5T2y99+pzzFglrAOJLXauGl9HMrgoz3Aj4L1BBjg48lVUj32nPUMg3
LYw7gb3CyE5KMeLuBzni45+oJBlQ2gpfdPSgLVNT+vIzGENT2cwDlWv02c+epzgt
QmClPNc/snwJH00LnGH/tpJcP02geXRDPlP2JdU6LNiTIZ8w6JgcP8cvhnOx7NMB
nuiUkxX9NLZc3jvA/O38Wm9c1FELCa2/NLMiM8yoihI3avfWS4hLUXkFbuM4lK8C
Nx2wfi7cPmmbV+qvP2SEgbgLb1iQhnGr0d6Ct5tv3rNeE/B1cJ3CJEL4cDJH2pW7
k9FrWz0OVBu19SUjyFWq9/KQEJ3SC8gIVO8IPJAZ6RvM67Nt4fTcdpa7LmWYqNsu
zVC8qtTsiP99lbAtJsXcSr2cqSJnBxO35z2t3991cp1KZJ6VEz9S3sn2wYlceqtu
270vrkUloi1q51l1Y8TF+kAGvS8PFDBUE4dVM4uvQqfjn5FIB+xxwJVRYGb3nE4M
p6Ocb0rPULhReQQkwNLupJDZa8nozUNn4xqji7pRJQh4UAIwW8zwTJuGiYjm+cX6
30cbEGmd623Gl1Bfuuvjg/acX9v/C0LKwCs65/7oj8CUliXAOSozsjFMZnmOu4wK
ask1uBvfCmUbL3YW/Fbu4lG4J3UpEETvutxtK/yolyzGbfI5ZtyTdFr+IqTbjwiw
Kvckmib8kVJFIXkp144dVsOoCalphjhsKWmc+hJ0QUf7IaKaLQv82D0yDJHMMU8b
OMh8CbVqjkzvppxeG0tVuX9RJePFtQ7GGYnc2IYgY2ifJitKIoXSQB3gPn+pVk66
Thcg1H4PymTIGbH+LPAnOgRj/V7SXsir2OE/tHfqrzvmzDsGtyCf5fh+8Xnbnow5
YlMrQ/oDvjQSchZaiNPiDNkrZmkpIxn8jJiJleHz5tTFaXhXJo1gEM/4b59itblo
HjuHZ5LAU6xKpCa5G+XCQlftrAZtdVROJ6GcJcXdubR/OGrEBi2u3eaRl/LHTj++
fAvkA9g6YdXqzzey9fLu1CG+48pqm2dBIPDGpFVnEZRkPbEtOODsn8/SbjMvENgp
F6bWpQ01PJasv5tKVMDV1YIlsbLgXEssBZ/pJ9RxerL+oeFmfC6Wm6uhmf7KEJxj
6BKktFVRqs0vkZPHkgXfmNcZz2zoT6kAeK+RuCbvvjS5AqpfG6dHiQCoMUOa/EMu
6x/vjm1stS/9OCqVG1QqEseaI1VXIDRUySZBSSqpdCwnWPmIQj0RQjPSPzsGUrp+
JdOrT8TTxjgUMbDygziBKK9QZ6dw/SgHCeAciXHy74iDsUq1uGiZZSGYExtGMHbo
BOqAoXLUeFFu4XxRUrqWfGPK65j9N3+8z8JgyTSxn4EJ9MMbu4lfnm40FUmltpiR
B4icmVdaRYRQnxtgSv/uz/eXyqBIHwvViebeU/e+RaokN0SPSvE91kF/hL01muET
PqenWdF6O3tvMPWKi3X2Txtkg/d/wc52kpEwlPOU0+907vSYUvXWS5sQe1gxCkS5
Y56YMbGEBttCsrRP+tmASaDZL/oP3pOaWcdAxOfB3TP7sVT5xz2ibQSixTvF/f7v
1/t0Di7N+ph5GYWQ3HBDZb1Ik9cGl7FX38jD/m0lvwQ/g+HxG9R+M5xzjxqh3dep
bys3KYx2DM3oXdFOm+eEupSmDtr3kK8VdLURDlOW/yKMW3GkHofkMoabKKlhF9BI
7qYbSSsEY2l6PB6XyZ5SVsI625V2YW4ZsYAjnMtfopZaBL3R+6rX1uVZo1FFI5QN
/2FZ1kbdR4vO8NN/DQS6fFXFSATh6KU/L3DZLa4E67Dpjrbt9OsoEANRC8jAuh7Y
RWWfSVD1nsBHzPyHdSrraN+ltADMnNnYc+3ZKFBnKFoU0tPYBdfDxN11j07t04wl
LlRfBOTW68GKwftDYvE0h1I9UvW1ddaT6AeJEqh/J57upVibdrzVwK2lld3HIUHR
WtZgh4FiLt8b3CtNUdsg3C1A+I7fR7ylWB+brmmz8NewJDDTT9B5I+2xcCL2IAau
jenDj6gbmTtHF6Ia0RDb/7bXXgKZ/MYLfSRmk+qLO4kePcNPOexuKVMBWHPNPV9d
HLulyBAsIuLq3JIY+Rylm4+TAoqxR4LHSQlFBGZ2b0uCXIrAn+YtalJ0viwpIw6R
04QRMn3YVo+fNw1k+NprXzhXzHv7U26oSYqgCdeW5Gt9jN/ViGUhsVgFlE2W4avn
e9qagn8KxRdPUl8ZKXLe+F2PUSZR49rpCfposO60psvWcDSznXOUnLid1q1CipOR
eM52u43Sw8F2Sk1ofNUOjSROAYVSfUaiASNs5VGnWNCSZW+U2YV01s710qtzLj6V
01NJBo/0FBfW0ZVqM51ubyb9Ufl4d1G4lTiMGSzRMF3j378+R7C0o7rw8uBVTCZO
yuI2/r43ChDzGRzDppoNrcVyhZKTxzvEVc7XTpS3XaiDBFYyJywv12TjA+1yKB8W
bFYFEG7CPgT68vY6Olqg6V8x2HfkzYNQwDMqbksyGJtFxfMYHuOXf1vqTchwtBMe
hWjt01SkPGDm3nGwJvWo+qWR2gfvDV5xrBBM9gimL3x30guvozBw9JsYduQxw2b9
3yh2d2APJS3DtDCXDWEYidkMwXiocKCq7QkWuiUyL3EsgxcrEuxZ2wiOhdeqj1XH
mqms+BEyUV6JUhUm8RhqpDTZEWMOZGw1I11CaNtKAz6qax9cxcTffZD91vl4TTNZ
/dpCMQAMAlF3FtdlHrjDoF3y8BdzC8WoMLmwjbXomjTC+XWBaZcCAO2wN2WtooQm
qejw1bFMUrjn4v8W/aAzVTs6ovp5idEdf6golwyW8TC/2EPIgoBXPVPEK4nNqD6R
sfDm4vAdnqEe5wzdaAEo3TuJyEsXI3JXS9DuYNg9RjAVJFN3ctwQwniIAj4ADRMY
ZKQAbXru+W2ygGxFZLmanK5K9Dl9oU1ve2/+81WD4NMkV4jQJihyKlcjdoIbet+w
g1jA/zDTMC4erMdET9ABL1u9jZ1gn6f6xV7Gk/6nrA6xEva58YlswZIMg6y2Od95
3xMEj5kfEAiZlTta7NuotYV9bKZ24jRGBpl1HngbNWLWRSFuWUZX5qhG/WhFx+bl
JWogPiWtoGw4dcpOkIxZ52ly6EitVznUzc07991E4YSERyH3uj3KDg/b6oA7b133
ROGiYyqiP7nr9zWWGoMT6K48e54Xb+/sct4HJq0LHRI8hjWFSGItPSqId7auy+Nu
iFRzk7XFbNHOk1RLSwO3ugyzyHvysPO9Cnk/AacBCWZRIckv1H0suQlTRHxiDna1
UaCttO0xGex69CmQBNN9TIKDUNLk59gIM00PpuBQKUqzK5TIHRt+4E0rMUJg9kdi
ro/QFO9Q2OOBNTDvHo9sEkmZz36vBxUgllaqWuH767GbYNoVqFJnNhjuoU+d5epN
/E0AIgSBDLhGLvCTRqr8rN5BRWeuBGAc6/8QKKxCSefZoHMo8n6KHVmViRUK3FZ8
ZmbfqTcnvmAYY1gFD114oR/cSqYjiDkAV6m0Oa18TV+fJiH9k6rk4gQSsmIeiypK
y2R2P/yars30mKJs2WAw3fhDk+uficrkpg6esjJgGW3tMtC+2a5ovGdTTfSpCJKw
N7xpMnnPp4Fpn3itlvuGbe93VSQK9FaA2wVZRKQC1Qrhe5l8YsMDoIgkWHSdvfKp
rzWv10vAXNAXw5x9gAWnK2o0RD+yvgqNVlaIj+zQIGb5tRwSbZSeEpt4LekJFuaw
+UnvWBgRYxSH6dSrvClRW5Qw/8jV4VneI8dJdmzzX4G2IQOPsthvQNlyeWaEYc5M
m8dacm6Fd8RZoP/pQogkSaq4X+ksNZpQ1PEeWCgmnsLWAAuS1D/ovz4lTbs2hitk
CO+r1nu82Ei133gzb3GwYQulutx9xaSbeLl9lLL0yKlq1PXI88Ai1uuv7tikzsPr
zrH0CqBurZ1QU4tcoeSffDz/f/LA1f+acJtzqHhE7ROljfoq+YleWWcJ5gfr2AxF
23J+D6BewREoQ8yVPl7UU0F7+8mV6T7WuGUk/MBpDsapF9grzF6PelIxxYgvRqSX
zXyb/c7ylKANZP+LonsHlLxYHLyqg4v30QH2pNvtVe6HeliPScOycIAydDmlgaI5
TGWZzpIdMFUWpcstEmIj3c1h7h5NKirrvCRnscCb7jW21jqx3tbcYt/6WAGBkBn4
XAFJivFAjUDK4znpB6qo1//G46a3ysrK5RYwqEuDNYRvK5PWlKlPK5Dh5zFdQTJl
ZDmD4CuNhIQeSdby/sWU5O+J3TIVXHnNqw+AETddaMLgnLTCDCjXBhZXrpSH5dFj
De9Qa3MpDO6ubbdC5SJtBGnTSCouY40BPuSYXQ5FvZ7CpNuyfGfwkDSiINSwF2vq
4qthaNYvBUvKpzDIdTeWnZOxKsaKez1lsA30u3TMjk+HMI1de0ASU4H1aqYVkxje
5zzOkCr2z+M106dGPj6/e4XeScU3NzwiGr9pQom47mV2T3b8331Tprczf7V9ETZV
SjpRCPP4Xg9Nh0jj0yG3rX3AokNTRs9QgzWKp/KlLyyF7NejinavpRAS2RZoYjmA
v/xsV9B6s5NQekqGTYlu6CsMD38zb15vaZJaHwTlqszC0botzYANBrMSzMc2uoEq
gEchwspdICvQKNbnVdr3De/ZokJr24Oq53t11I1zEP95T/XFlAAWtqUptBpvrxRa
i/3M+E6MRK+KR1EguVyYZ3bfBTXLbTYD3QyZJEKmQB3MkaL1nz3D/bNHYKdFiCes
wJwVyKWjp9MKuHTgtoGHqLsuqIWjydoERXQYgUIFkCcNboverj6rBCL2vL5bOiuq
pQCkTagP9yZdzWGzC9KTx0NpN2y5oP6bRVvO7o6I06vBwxstwukpRQMrVbN8Z66G
oNWrablL6DjATGUTO6sGyrcfDqRUQhMcoZBvuKwLqIShAolB2rkoz0uMXF9IFRd+
qFydnqUM/t4wEnFcTpERI8Oy2XUPAbPURh2Zm7Kd6hQNwGshslD/TEvnqTFQiTYK
pgOaaJpGRHCBKxLExRYX60jmKIO9zzD7AMslVhHrFIsuEb6rV0hwK4MHw2MNReB0
IXvucbu+9mx/Ql6L7l62jnT4wgiNt8taCPlFeW7B8QKqQBfL6yEPyO78Iv4MRqqH
wax8d3AdTK0Q8bTT8QHJb6cedvQbiLnFWky5K6Ygr4BilC+InlFfMgMSxBVJ0YqJ
hYn3g89rr2XCf2yd6mRTMenJSL3EFGZZlARs+31aC695J3QsiudEr4KAMAuRJgfO
qrZYgzQG4iv6A/0bNonqzhf25Vu/y7nsokc8aj8Bd2mw1vK9ZSXU9100jJDDm25R
AgKZL1HbN2FcDYrgFFRy3dDnJQrA5ktzetvDMd1w7z5mDIH8oUtPr8b+ZHdtEKgW
wB2W0RYo90CRB9P4FgFzz7lrd1hbTJBG4T4aTlJbvm8618cc6mfAz9uYm4/zehoN
SL6xOXdQfyeTihMRS3OTUVjbzFi6u3pKaIeM6+pPkATf0V2Z831Ub/eL44r4862c
Z2JInxcyWaKb9yFHdBUNd/szTI8Cb8El3VL8TNLddCfJ1uF8TJtxlZ23nuBEY5x2
4AzJoGEkcQNdCwtburWwT8FUsegRLIj/MbzGOoYQ7F4Vn/vhweCdWdtwHlsbHuIH
V1+shbGrOV288jEGL4+rZKtOJh9GP2lQFozCuASRb+VzR2xkmeodtzqYfXNfbzd6
hRHJesj9UdnF4ukf40qVFw9zaVlo85pDizx/e9yxY9z4WzcR2kF3HfZrR/J18I+X
xiFLjYq4Ik63yHJK1NXo+tU3TY06AsrpIO5yvgmJO+5gw4TMCxwmlQchS86nvUTz
1x/p06E5ntUzvaI0unYVZe3ZwiXmDTgkV3bjdAN/R3CC1B0W1btnxUyuJ9bFsaok
xmZtddSaSR6c6Cl/d5sEEiy9urOIN3NNWhXL7bJCvs5FcmfvNjJLnJs2/d9boAxm
3C/dyii9/VdqA+aNBYR9m3eLltkKB0XuLhsVfc/DkgwGme3SZZ6+IHTw27CPCJL8
SHzOEKVmVI/0e/s4EZEtsSsh44+IzuZiNmm3s2h+mE3tOKFRt7ZVaXTzDI/QUYxZ
25YpkUXVNODi+Ywe5LgJWwmNGsEPxFd1wagU5i9X/wglheRThIwmNUjGv0S4jDnP
QyTNsxgcI+icnK8VLrDlwS0Za5q83dDxsXLUtWqbG9ME2GA9G8q2BEh6oN5JqVyR
K1XIKdJcy+APEMZNMyruYecCPnonVtP6Xx8Lv376Bkup7W0OZEP43CwQPCO1ujyS
JHaDGrmmMTSi5sfoXIPi8dTISbjNG9KZqjQumFsuBAzIKWWfVDVwmiMe1zOI4omf
uql8WsYLftHwhr4sq1Y4TCMB9aUCXlgOsd0pEylsh+ybugfzMpecQBWAQuDOBAsh
7D1zL9/qERGq20VZrczgNk74jwBIhjTp2EPjxEY+dr2Zokp77cDivTctfLUHeJke
tyqjHQFLMVcNR9d0B//OM0BSgKedSQVbFGxPO5QWqCl3IdbAqBWEyuPpXWR3fL3l
T4O9MgR3DtrW24P5eQ47NwGLA1bR+qWwz7S5PbJ3Ych96PbU/N1Hu4R2IXcqM4sp
4IPrNDLY8XHXYN5ox570qAVgYZ55pbcXHzRdIthq4IiX3mMVYCZwjSD8tqwFcFlC
jA0H06g0gK9lh85VCxEYrSRw+2oHOAxo9cPWuVBswVwdb8akRWso5swDp+HP7BF+
w/FzUGZYghxEBGMTQ1LgfM58mglGvi6WwlsaTu9Iho3t6g6CK+aOjUfHSL2xWBhp
Wdb2Wwn28f8dJOlPzDL7YT//nrN/lCAWeRU3E5LoqkjuX6PkzBtiOJQxajsGcXLV
/qG1KV3pXJm8/XkRdVuxgVPLZ3Jx4VAfa6MkNvEVKfZdnqaHaCtmT5H5LBekT/KR
IaYeG/WWMu8hT0ACmOD3cNeJhy4kFBcRThIHc0Piyh2zRcVHtGrzqfF8BXfTzGTf
/C67+nyEC//1Vsix7De29BChqsWGBcarkUtGNCTsJPfh0ETXh/83mKgh70s9vqzu
XNg/4FOp56gl3Jv5sm35o8SprvoUbkQ19SWaxs4omLQXVfOJ+aNqC2J4eAqY+9gw
P7e8XULa4pasBBbU1UWlPV32h4/oSDbrJa1lTCGi3gyeYUp6P6NtfWHfX50G9uTD
gLo889VP+4B6vE8vPuP+GpEransUYpkgPAdaeMBuw7d1oueye7xBs+zLBOBBsdNG
xEKfcjuyrKK5+0p0cfQPAjoBoBfBLNW+m/TWAmYwjrxI3xPAXw7oblZTTHKK7H2B
RPWS7m80c7zugo6mdDMm1SagArg/VIk73aUI6F0mHJBBCyLFpF3VAPQe3SDXSO08
nVTmDg4xoykUII07Kinn519iyPb1TIUvIyRLw6z4TKGWLjS2aC2+1FP7YBNOiaOj
cS12K4yfEEUAelZL2XdFvvunT4Xl+cc1pcjspdg7mlw/jLjhZ1rcjHwmjui+6fz4
a7F0eEt/XC43iW5eoe7ASYvm+iYPfFa+A1NCFYmj3Da7VfFYRfKrD9W/YfjcWorB
X6bzIQrD18Xu8/TGOwjFp7IWwlWnb+XBMNKRi8AnzQkNpjOPVpxxua38BUkHX5Ey
RVm+w5mcAoEExFRQgMNo3Ipg++av1epYxGUCC5x8qIO1r7dlW/WPkimOVf3el/MA
M1bUggqi126SQvnpuSr5IJaZqs9ihhzoYcCImH/cHuGjJe4BIciTmNatoLU55v2F
bFcmcotPp7M2cQ6ps0bzf0RvorBP8GXy9OKzbjPElzF6J7oTuhrVhdhGos1XgG8T
DXpujeOJzQcVUayCQ8FrmkZHGoZy4Y2rZ4fh64Vy8dVYccq0ibjhvfMdeMx/Fump
5FHLU8YwR9YIaSyEERi1G9LKmNVT5QYc//vwTBM4Wx7e6RDqj4qopwgO53+lhb1U
mCMU+h7Ivaxr/Bg/77CQok9vvzGBHk4zZsPQcdNdcJ+BLBnyjO4DkWUpsG31jH2G
UuPYWJAXOzwNFqvB1ZuzbJxIvzh3YpxdehiMGOFOp9g5PE1aZEyYEf29FKCXZjSw
Ls4PWgghKN86kld5Dal7JWCzDwfXCuyYafLS0SueSuA0l+zA0WS2h/Eai7uTEgC+
enlM/kOdeVfMmP+S/07xPNYDgHB7Y35Kv03x0WVjZGxtuYhEsbzS9MoUXaachzKs
5dGABbQ5rIiBxKllDQjqKLpc0aYrSzjcajslH7wZelWgc1tKcYbhgjI87nbSv/nB
MZUUVCGyLa+bWzwClVrgpHfFLWlR6E30zmEeYbvppayXJX1nB0nKgsUMzoxHkmjF
fy2LaCR542t8X5noT5EV4YEsCXwcsN4VPrvJ7Xmso4pAyT8GdIR4/6CfP+poIdCo
sX1ku6spDqJ7fUimbOIr5vqid+8wsiJHUnWkU4jH7s9iCIrkOyNruIQukhiSdgpe
6aIzMHRo8FtkGnh8e7sRVMDQKsBeGgf6xHUILRPR9FWpJeAuvTrjRSp1DBeLvPgZ
B+vVvgq7Id8lmAzAHTaFASWviu59e7fNAJJzlVuvRIsOup1LXnRxKxR3C6laHdTY
jpuF2xuYDQvRyiPcS9xOXKcWsb3AGWvgFmoJCIoZUHDOoj7pAYgu2kz1lpPZqS+E
xxGYBYdr5VL0hYLFVc05ms2QiKLKnAjw+3GDWgrR+eNKEoQKcN73jkSp0tOCk53r
ySypXWCy0opnZsjlfPPQL2OUilmsjXBENlR1LZY9FGAJItHFDilKHDEGda7RDNLX
QPw7ukV3QCvCp1UMJQuCuZe7DO91LUyT9XX56Vhv1450/uxho39FpYTjAc8Z8BDI
xUHZGkYVgVl9EHc/qBm4wW7cKVV5wqktQqsQ0sg7dLVT+s9q8hMeWccpqAzvwd11
g2/1nKNt00j9A5i3AOD0TOjWtxZylAthEVkUQDYYJwSw3OGelMtKDxwpSy2obA1z
R9UfZ0Gq0cU8MUhX5+Vjz+088Wf3p2JJH1HSknRDoY/10Qcf7NJ1ZODEVJk+pgYF
lRktG+IPrnugrXUixp4lj7ZfbXLTJRUjRpDnRltwZHloMxOr1rLJs45F8UaJuLMF
1+PYZXZ3c/tZAesUJGapyCmHfKSLDXw1Gx+Xa1s9qzEaM59myWIHt7jdoym2OkTJ
IcKMSkSQ07Or9ApNB4LW5KkHrjrUBDsgnrIlxq4PxKro299vpzDuuXzRZPsVJcch
lWNKZrtPL0BEzCJyLJ61zXQO+N7qnUa+sEJIkh35U3Rebr3TV6ci8oWOQwCpEbBU
uLs/O9jh/XgvKIChnkQs6jU602rSnp9rtE/UWwoUBwTppgr5j6pAY/F2GaZ+T35T
Tk/xWoIUy21exx2e2Is/WjiHXrYLhQ718PgU85CeXeiMrzxU4ba/rWFnR/57SqRD
nIoe5rzWBlFDG+ly5FhcrmsfwCDlsInYKtNxvDiDaxuCtfjvNYZSbhecGdcMMPBB
daxj4R42siI4FIlHTl7wtiAYQVas6Xh3g2FdRswSJ6p/+pOCbVYPZti2/aGcBRcz
iTkTsfaQJSaLksB3mz7iCIbMJcBPP75jxErkjw90+C+pruQhFeBTKKOhLfTHKChI
sGvjNcIG/9g/124P88p04rQypqf3tdXAk5SLAEXHlT1Sg9v3HTMrMNbrit9Wm78J
A/EMd4IqnoEez3fiIuvEP88gzg71PW6x/Wb3CaXfTEJTyORVwoHz9IxV0bSc5pbP
8rHsI+7Z/yw83vM3XvxKNFO/64Dox0Rc9gHcX61eraivb6L8yb4UeTtVlIViGzNz
mHJT2oOQbt5RwIxsfpKKEam1QkIx3DL6LdGTXHftLnVVO9Ad3/82qy3bSo5Svqb9
+84X6fQQ7Sg2lzrif6sTryRHIAdjj8kRP7zgn+xi2bI+dia1bMPWhoAUSQaLVI80
JYermGE8MJX09ls3Lo8kyHpcanfsAoFRwZFrVjFlam2LUwxAaikGV94KLRlqe0rx
CCB7COlwFY0Dbqvd9Xhze1aFr+yXP9NAnoenFtqW+NbuvBB67tLHvIeJCbE9jtkK
t6gVlw7MPCZYFHN2bmZooBIQGCXL8QlWxR+5lncALITv4Zb+loCUUOsRJ+RV2z4Q
jyg/bkWBzbQB0hLmE943sO60E4OHofp9OXnffJC04phqgHk0cZPvK/gX5qiM/O5d
54VvyxK3SkYihYXcK5dcgd+wINjcdLzIsbEpW5DCZPne+Y5P7dV8afBt3WuColup
Oz9qlHgFZ5ggdjgcETPwhBAJ3GYDl9OkZUFyf8qG/DsyewZSnI9qRUfGk8uPadFE
E+RQxLbBVlJ5H3JQd5o6lQUxNjy7E6p19RdSX9nXSOn6KxfdljzaCxuVn+VizsaB
40rRPHugOPIXa05euTKYTbM69sHnPfV2SG9BM+SmLVTfaLaPWT7+jUJHZPCeaoXy
0Csh83T2SEQxDwreUPhtMbUaPq9YjCG2cXimf7Aol1RCRncCnYVsznojWkpN/s+L
7flna9gFobmaj/aYuu4PUCG17jPfbfqmZ96YLo1pbNaYuHHiZZyljnIr/nqGGnof
BUJ67YqbWhKY2xbC0wz39anurRSlisgTvXNu9EUFYQMW69i+hrOsDqjVVmWfGZUx
5bB3Buu33bEDin9i55/cAcOqTztla4x6LyRuSTLvAICz7D5t3jJVYldl8B9+kMeu
mvn+REQNYjgpSDzWfwnxqV4qcw1EaHTU+plM3i3CFQBA40brr5PFpEJtzORHADZ5
a3wD7WPvABsxIKlXftVg4Y5TrW8kVK3m/5uSvv7DZ5+5CK7bK7FndbDvNHQ3qQkf
NaDDFOSghC2etN3bPLApPMLbL3YNat8M/h0Z39oQnL2cgElvhvfmOg2wvpTvJChW
c8DDxERy0dfMcTsoL0bpI78i/fcXOL3Ihu3R4n+2mDvcbV4fEUfi2qiX+JuqovAB
UcOqKz4SwG0RcDIZ2NE1+mQNfjia+aKqSjs2pIOoz8ZAFpFEOCbHtoZQspsAetUi
ID/Ai+5/zLDPaoRL7B1kjiShOG/9ZvB2+zX0q3i249pvsnGhv1xNfQBZodqYN2Rg
MQKO1ujJQSrpk+OiZMB+oS7/llmKo/mDSPRQVJovG5aUI2bEu8A8yTVXQYmr7Ptg
8BBNAwU+EBcoytQTPYwkhHuWb0z24eQHF9q+LDoXJHeRNeDOl+MjqWwgsrYvbDBO
oSOtfiFWUhPjpA1k36fyiYl75uN7nGRr99a9hB1n64jVAMnedjAV1Bgchyj7jGiu
uTfgxHOxs63gtWZsNVjZo6erxVO9M2QL08MHXY5DN1aV/MUADkFzFIk9tgkiCpNl
k4RMO2hhd461K6fUlcGQ+NO24GImFMlC37rPadXCLkLgB4K1KG+gWuO2bp7l5T/6
c/ELzgqvMKuZg1b++BPI+Sg0BFpb9HQWs7Vs5KWXpEJJjWmGeqfyx6KYJSRvM+7q
NjH0CSPEQ4LoYJkI60xGD26niVk4b5iCjUZnfu0TbnOPLvr0tlxdCsqNXPffVmHd
juCacWFmuSrJ95VoX4oUDP56XcnvEYIWgRGzIQNbo1A7LUnpv0yMM5c3g/g4S+KA
FRqAJoeIdfPw9im0n/AOZfgGTLY3vWDiPKfETLBNZnXP9UTsYlWf4rqIFdcTdJnu
qznfBA1Vz1oSnFX+dY8ocImTEW4BELnDwtwqY1keB9Mody3jYROO5HTPQgbuobpn
ZVI7y8xkg6xR/4rmQ1BjWvOAF/eP8/oH1vn4/GYGT0Fk+2b5zXAq5ypIv5WoSGAO
YajFMJLwndRNHYdAAMoDG3T/ssG/3ZNspFA1d7oDuWiOc41zbbamF2f8u+YBBQ7U
eRAXNyqrpJGtOYtEb8KPAmumdKTCLEWaVt0Fm+d8O8Lqqqmg4OvYHaORQpLiBHSp
pGEyObn9y1dn9Bhyw5nVtPFQBDCn9h2XAIa+ZgeyXsh+GOyntpoTDquMCXHHI6NQ
49afFWzIbjAK/1YetxVEl8Zp88/CuKrWNR0LQPBe1+2yVQi5EYxIgHODVTtQeSdB
dGqkO3Fzc8jnB+qHJiFBU7AoIhJ+8QHt+3VILN4f5fA5hddlAiiH0HEWO9cKIkwC
pEd4oYP7iqhOh/4DIbavH+UFc6poVUcH+cDSU1BA3Kz3H+k/FVCM4qLO6dbKyQan
8X97lU3Yt5OcWNAUlkoz5IXMpRzJ7GnWSW90t0MDeQYvOR2HqZuvNuceyOCBkkFy
sgp8UdKfVkPbC7Sv6781/7ZqeERKAS+bK63Br96kPfOl9I8SFaGwKYWcvzGtWLaM
xiTkGU0xLgYKg+n7zKGYsBA0W2NTzcfMxg5x7TNMoNk/qzuKKULEs1BJfqdsNNi3
kN8GbnGFTc+elg1XyW5Vm4ZyUOa6pY6/LUUEs1Yp/CS2SqeIpJLuUXTRD+6RdvCO
VIokMw12fHPU20dO3qp8CGURKmP3NCIGQqsGtMLJR5/f1Ke+/V7U+wuIKSXAPuWA
hHpA+WnHAX3Ju49LlikZ4kQH0LQ/c5GSMBnrajmsu7p2MLdliAOuqEdr3Own5A+1
dgC00JjWlFSyHmsjFOBtGI+f2pXZwknLgVQfZS1j9kpfFWxhParGKOrvayeg3MfF
K4llTfnNvoNJs+FR5Niu+uZ8m652EWXCSikDWgSKyGf5p4ZXHvNM5CKe9ei8vVoN
byc5cqmPQ6w9sJAWzsvisb8eKqDXQvCblwAybgV7xIjpiBi1COER6152jnGT7hKM
zEE8S3HsmqYdlYFmIaBrSHuufXHj9WaYF9QoWgLBA6rbhW8PTsB963kWhNiY2Vcy
HY2NIiE8iWm1FIAxZNXsVGxSBmdpwMV/H57J23TTQBFN+ox407fdQrRaEU5+gGnk
7HNr1hbykjphPt5EC5se3NSzl6/bis9z4y1qtOUQMRUAMSve7YJjphq5ySYVkLXv
gL7ngAot1bjopnjMoAr1j/Hnt59YXWryrXfGmUnvDqSS9Se5fTWBYRfCrWX/CJOA
cG0oXgMKUDRVuuGg73JMTJmzu1XkLaolvR8DAD+D6hFmiJToNdGc/acl4W2t5IZ6
EmYPV1zWa0kqLMZrIkoqOTTMfG2IXviygy4FxLuJssd+CWZApHDDVA+YAbmas/80
ZFJt9j3KlzZHm0kzqJKnQwzMPUKP2o9I/XW2er9vdIn/jX7X0s2cq7nrCy7DUf+M
4kgBWFgPQLPy1oDgCYlGriEwwAV7/znieldQo/Dyywiiy32zkKJdoNoNfHJN3TxI
YRKLnCCBkfpSYBdfR239R0BsYXzj7IxIowxRVAGz8phjcg8PztdwWZ+uB4/nMMsU
zhT7qyKn7auqXJ8N+ot6h8371oXRjlI4VRWBzXoumnCazBMoEWE/NIKBtPBE6XE+
iLsABzHbqbb5S1BPb3Hw/ichX8Z+AiU0dOZ1qzW31h2Xi0AVNd9gnAWZHM7EEa+v
6Y+WcgXEMg2kBj4EvH2HCOyvvlcPoWver0ZDNQDkOw8bOOxWMWzes8rd6HZVfAvI
5zbuEeck5hdd5m4NhvJM/whCLLsAcmI/yfQGEPvVl18PbIZ8pyvzLJX5HqEcaY5U
pW4wCEBeXQYFb88yt0qHXzTX3zAFYOVb/Ib+rOfVrLZvxNECxxWG/vwUkm/KaqFZ
Nq6+rQTD9SrGLLlv2bbnEzyH3D5cqtI7tqMaAvRpnW0HMWRl/F59Bhv8m89Eu5v6
65SVm5BLXoSKh0XUChJ0Zkzi/vTwe7ytAS6KouaxyLeO8yARPUEds/6rn/nKBDuo
i9hZydhM8xkowbd0p9ou1PhKaZlXssXpHvl3edUkHiCEhNW/2uuPIbYUykMm53gQ
rJCu3G1Sc1jvphGjkTSSN/qxEYPWUWrPSZWZoYVxRYRMc8ictaQ9Y/yC/iOnxjR5
w4Ogjq7MdduuM2RnS5rrk7nPmuNsVIB9q4XJgWEVkN/eBRyJn8ie5PAgYmLT0xLd
ylSFRQfUgtK58DqVFTpnP6hDgIZCroP4qCw80ZakLn6ZiGN3D/Fc4mQA8vyNIq8K
SN0bPhJ2xN0D82j/kRumWhmoPk7mYiDRXBSxoIE7Sg4FXJohoZeNOs4t9X1b31X8
G1SQN7CNWDQTLBhHP+GawN99IAamok2xduExcfn7mDuDpl64wgj7hgtVT5oPje+V
I2yYBIBmmZAjyPLKYwsqSTt9QCzWwbKEZO2zIVBfpM8G17suvuMo6Q88z3axvtMq
7jJ3pTYngji/v5WcdW5yL7fR7DcbJ9EEWE1edNf1UOOUda+j9Omsrz9tY32eNL3S
EmOOWyMQ0GItx6ncFf2jv8SkVo3gXO+4M0y9m2S/hSsncd/nyX7rBtd2PQlkJqlJ
ZVKrp1lD8sDfl/tHobRswUwT9hV2UGTsGqmq1hiSoPwI906eKGqMTseqDzid5wjX
OfYCWbgMR6TOBNULY3TEMjnXsiIEljTE44sbs0XeF6qho2jv0vKj6UUUWsBQ8Xno
KOM5nJHG3UHvdVOmW+NsqBXPX1rAUoCrTZzdCHkp6wYg6ROJ7sB4v917Sk5NPkji
6efkxqWWkSAkQto9NYEl++1kP5R1M37RlgGwspDe1Op8s5dP1LXl1bu5ak3Dd8Fu
pRctwV7S1IAwVt9J+CenU8HPlytZzpPF2dHiMlX9ZSBQkYURmbD69GnM+ANtNz8H
7l47IaWgW0LsqGYy/9WfosXaRysv1ZFJr0Ox46A/ynJABHOyYC6AuD3lz/tcTWpt
qQfjBUXTeALCJkidT+gpGETE9vOzwz3liclLPekomCgEmxUF7skkcpVvjArQCFNs
SWdsEKr978n0Q4IF68WJBHZSSjVo/a+I9uRJ+Q3hxZDRS17nXvVv2rliz6p+pKaY
THFvNUtWBfB8RyUT1tR5qyvBGQQEhsgHtL2BQcjvjWQ7i3ABmQo5/Asc7TTFwyfg
YIRx2WAOMooVH30ZvDZQ0Q000cd6LM60gtwdBG+8CdFxocwr/qZSWX8gZPgxIra+
JefnCYPlVGcsZY4yHHHeGkb3Efh7qzcATI9PeU0bIMjLF7yNGmCaEngXVQ+/cnxT
jiFfA4WEzCSEfend3C2NaqJFa133v/tZhQLUEJ93Xds5Ec4V6Yi2r+3Sxr19JjA6
NaqB5Iso3p95bGU6L4of0bLjCOs/aeN8kmGItEXMBNMYuOCWz18iOgMldMm1mYXW
GrGWJrgCP2HMNPWvOX9FJgFY37b58cn7dA0hC+fYA9CKvDpI1jrqVysIII2Dbs6k
eSHQyuVkC5BQOaxXR3J7KMYdrJ23CwrLU64sgdNXd1cGSi61boE2+SKNZRvSYwNo
FL8i+0JucOdthaTTzsHuxqbthyd3xUaMKi/tzvhZ31SwhQGbVrxhUIYaxgleFsrE
VUIAuBeRAoC2Gcpjj9V7JhASBcmq6o/2ukdzUlb2F4gga8gUxQK11WdsjrP5qu9f
flaIQLtuJ7v3gL871ALNwoT/tIM9Tjof8zN1y1a/HvfJMqLUbfbHONVFzPDkGFEH
5Ak8WTrt9WEF31mlzMfZLdh54aXf4hakclqDgcJCrXdbyC6x3cOu+9J0sQkS5bQF
z0c41lgJAj1yCeu+YR6c/0inTX1ry9aP7WNGY59PtvPIZQZGlvFKH2mf2sr75KDm
P6RVEOnL+p4uagNkiaqCloOgcTKqMNh1hL72NIPqGqE5EPCCvk/Fy0+p/+elQYPx
dXfNb7fyfU3F2ej1kyvuT/9z+6M8qbxgNy5Qihv575a3Yu/6Ij9yS7gb9oi+Cn2F
CY7ehKPKKs+1EjVoA0uogD1T/fqTPAFmHFu5QqYUzJWHsiNK6tHLojO7eVccbbNh
spnQCw0BOeb3JXgFYK7OaEyBwhMwTNP2ggPFWuL6V8+iZLmNjniFBgJIAs2SFLhZ
XLP5aEyaIvNOnTjnJ7/eWvqojk1FQN9slYql43idw9yLKTWldxxiIffw5umnAZt8
rUj/VVLHGy3ZJenFvLJDR57QlRcYw3ocuChJTCjb6sDhIOXt8Sfl4t3A+AdC3Tzq
1Xk6ynSZ2lJhFUK5ahQbwBH0g+sd4SkxXB24BxpbIcA5YAuO9Opcmbqj5AzhNDS0
M1DFsL0d9F+SZJx1otMWtqFE3H1nYb6c4kug1gkLtboRnIjJ8ujT7AjUIqGvbd9i
Tx0MywVEAE/ITkT2iBwGZ3Zx0309mmkHN1445AEDLrkbxqfb811aRCniSeIaWqGJ
eNKp5XnYLXBFOTirLqcvS1iKH/arvHw+5uhBPIY3D7H0HWewSzLk/GfYISruSPgL
Mmb1+WVG9asolDwwJ1Ksk0kLtnPrIzKWz6/0SEvEMzuBwVtxhheWSjyspgVcWvyX
w/8dUrqQwm23yQoDrE4G4bSy7YuMVHlQndLo5ccCAvKF+IFFj6+D/RQ+Z0IjmH5o
IOWbs0i22aEbglfGj9C2uo8GfMoRtCDUK9D03HBGjGbvvqV3sISKjzqV5AMnEHYX
GCi0XSSmCG1DKTt7AC1XNWtnmeX73R1QPSSlHJ4NqwJOJHNjiVZ/5xYsocbe10wQ
aEqq8nTpa5Sa4btQfzoMvH6ez1d7BtTHezW0wp0fw20Nk1ZPZkBuKdDxq+ZnOK55
JodEA097NGjfCuU1iz52uhouRVJmFQDLXmP3sXdYIOJMCV/KR26OBLljaGqO4W/G
uSgHm1fqW6uq1wwMVdkOPts5prbEe3ftwiRegk9h3CZAzlv5rgxinRWzDZ1vD/cm
W1130c1jTAIvB8hWInc8CDStl+TZ8vrGsSi6GPc2HmJ4L01c5tmkc2zxek5ykw4y
GPAp4SilUJ0WxTEdjz2NVvEH+A4hLmIibYa2IjtMl3SHSKxkBtb/qa6Su1IDye4B
Qsh44Y4mGVSFmGUyaGj52FqmPj9OftfGS1gYu+JdJPNKyrbN8iKwXWl6SdBP+XfW
4SOyik/7Vr+OjBIT5mLZmbLu8/MLVSGqrC35hLwNTG99WSyJVf8C7dPFTpNSTrVh
pDsADmNQ8DVUriVpFbmrigUklXO72XXFtK0yFzx1HYWMfvOhxfEE+Q1PJQQFZvoT
BCWKpEHh9O40fyq1mzRwmJyX7aqVueFYphbBciFLedTGG6myA+f5wj+qX6r3TBZK
ei5rqEIjQ8PDajfdWQYj2kcRC75P/cabSoWcRn7S3jHM55p8x3cUC4CPYfoUNOF/
rsMlj8tMKsV9zgIao8LCCelyCbiKU6RWV06FLaf+ebM4AaRnMWsSLq64LVGG/4IK
E6eFaThwYWefT/UsXF5CSAnhcxM5zYEX3vhx+SO0U/5P98BxqQ1WqkRcJzL5yNM3
9lvmkTg4BgIC1yC9iiJrZO8Fa+n4MbDGG9vfnj3nnzXbtlUZeyF25yXpl3c3vl8P
b6cZAihwvgi5gAqAE16A38/8FKhsLnUBX4k+v2XG0fHpQAQEu28wR4zZtNd3jI6b
4DlFfKBFnK2L0o4lTymGOWg2v/vHHj0C+G1pqRZmWYYnD5zK2gW5SINfdBI0B2yx
ENKowAw0RnOq1lWWcMG7XLxFEltZexcWMJlnCi5l4CCZmwquRRSakjbtQExxzb3Q
H+e+oPowNLBVAlprD3JkOxPaABvs5oZvMQW4A8oDCjc4WahFgi6+NHJiYdeEe7v0
WDuzl4lucXMeikln5hi3lHgJSr+eOspsNxn8nV8/P4UOd99JSV/PK5gd/9felZ9C
/ufXzCmI9eQCH90XG57EbbSEOa09dfbKTQiaqSJ/CrznKNhwdTaeqTC4oxWEHQ2Z
luptvG5cAP598ckmvS0ohgpWhMk3nDSqu8d8iPL9OJqj7LACkI0deGdzwZkswEjD
f+/JPqalYR9apHytkNo1ZVG7zEx1y/X6Lv502tPDX9GvDJ0LJodRi/KyCDnIuudZ
7hmcuLvspHnwvUrlqIdovQUZ3m3niYJ5Zknv1dx0LpTxVAAzSgc53yIv3NIKYXHW
3lKpnpx8jToqZDRHl80v6/qxp6ePfXhwTvo2o9/m1kQegqSRxbZnSr3SyqPB2P4a
XY19f/xthKED8jy750ooFfL2/JquvhikzWR/kRk1iuajP24myGAL9GHQSSLohykh
643yQXRG9JI6vVeIWWgdLUQnR5aSQgQeCQECZmFGuACFqmMsh3Ov1P3VvH+Njhvz
xsyK6tJm57J6gGvKiMgBzJSvQODlK5JJV8ahSqSuaxcK3FWP4GGskBdRjGaHh8ao
ZpW0QXSBGYEt7GbSGlUbzKKqsm6YO9+qLejeM69AkbLdkjhnTnsK5M9w2RZmQb2o
bGXIzSwglPzNL+Pd94CXyEmRFJGk6+twmZof72cY2swcCYDTZeqn8w/h/Y3IhgGP
jhchaAKOZqq3Pgp2TSGMZ99pya878Z4OL142eKXeal2cHEW1j2gpmNzG4NrtRE9K
Z9rGZbdmhmErQuddEwh2RGgnmiCGMDK6Krvk6ds/qGpqMvZM6Onsp4WXKybkotV1
+u0vzaezlzjoXg+zwq+nFuif8DBj3c87CmZx8MYnFwOGtwaQqvnCYiWmoxpX6HWu
thAJ7aTfDrw6p5JG5McoIe2q8e+87TkEjTtb6Rj/Rps3opcVgX1bOwHJNEkPHxLh
4yBKdJXwQHRbv3YCCMaaeC4YubTpMmDWqIR74QzS3Kdi3/Abk52ioZQhRYwCi+az
+5nP9t5kD51FmzTJp4PGUMIeXPzlIrAiatNaeSrvXfJzeVW0cAU9qOMCAdxD4dip
KdqQ2EKatWOR1JJmWUC4vQebj6vbMsy6XETeq5+R2EqI0WdKgHY7k+AUrz2p1pa4
r2luCY2jkxn4rYusckm1iiaiX8HDdGvnRqU8pBR6oLX8j5CBzB/KtwKHnoyJDUCT
Z24LmzaaYRUjkocoowdMOlJtcTITPXSp6ej5d/hwkAdwnKx0bMh/a1Pygcd/8gfk
UcmFVZtPP0bD8SoOLcefcysoa4ozWXYLpYYeVBxJAVW8St7Pmgaj9YB9l2l4NnfF
GT+0SaYAMcGKDkaMDLqrgBtBIDbKPLmCmdzt7Pkky2IABQvk7rhktu4a+O7K7JX9
90B+RO64aTaxKf5dWYi4sHMQxGNIlNF7ScGO+2jsWXqo4mYrQxgjrFWX9vqsKLuD
JYQl+vAZBMTFmUCFihe/H3/zBOD79QV/2wVBahiU0uqnPLMbdPjHk4JKhVOwgK8/
hf3e/csjD5UMYVXf6LSxJsv61ZElJitF/s7z9Hb3A3AGVRBN98LOZWPzcUHafxA0
uA7Dc2Mk/flPB/V7WSvXDhxjLWJi5KV1y1qKcJQ716dSKBgL86/D+HIRqbQ5nPvW
A/senpIi6/G1GzIdwTEKWUfjUv5KoDXAQos+l8rWxJN/a4uQMnT/Se17/k0F6EsJ
ZfDnDRVTVAhcruasg/H2LlESlsR3B5VE4aazFQ59qy36wmJapFVlOuzylc+1tM1c
n/DoKsfHmIvbJ4+/yxAt7HEukgnObZQjORpWEwvW/tOWUVjl6U8ZUn0/uWON32xB
OV/LxLcfYflgMAzDfjyyKkROQ85upVkwmm0fPednAQbzSfH9DQXp8J32dS61vcth
Lt0VufDWYoNwSkywI/ygBqCV96Q3neyjPaw5AerrzmeLgRvCXqObTRX8KZlNnMz8
NgBXtGB+7pzkbVlw86+O+EI2LH1MO1LAJo0FsgA6WVU8iyeE+RHK3Y3AK2yoX2Nn
D/BYGcjaVJQ18RV+rQEY46LMP2lsbOi5KuJdhbmQKnAeTWaqbxR45S7PGwXKyj4V
L0VC70Mojks8fjXRv1uE8wV/PwN0iqX3V71+rwt6mcKRBFbh7mKwTBBDx6uTeKeS
ZIMSArMR4qTEhl1+Xa/6kJXo4dW1bQLMA0/KGELoIoB3pm+g2vXuV/W1fLXSdvQO
6bu+bE0CCQddQ0IX/z2NtORGJWYGwTntmjd3iEfJbLLoxPiOdI2WkQd3aEAzH5vr
S+dy92Jxo8OZB3ufFN+JgVw4/7PCBNF6wJuhpr2HLmA6mWlvSZnkYU2QBgFgDFrd
jWlVOwqmt4ZeEMqWd16KTAUP+dLoOxNXL/5aBKCLXZYcvGz3+8auekfnc5aoRs9r
WAILnQmijojNTgJTPocvblXDK1ESeWIbx0rCAXZYtDXqRAPAwadiSBaIAkunJbPJ
avefgftgUtj0roWWu2k20WSgGAdLCQhliNcw5vfSyGr3+4MtvbUUJiCA3XCSzGQ8
LeUmwehwqqeY6X+qcvIay1plAY9mkormh/FLxTH2NUeFMYHc1EHAAuCef3u9kLUb
Jm4HMCs8qoDFtlXib9UL02MiUNP0yEcGEgwvGWIq2PKOUQJylvAX5huXv5vCywws
GwujWZFI3tqwYkISe9xGjPRlOPo5H5WeZKmvSiVoxziAsw+dM08X5fhpX8WN7Qbt
Rbbk/Zbya8Ym6RYpRSaQ8MWK34qZuUQ8oqmCSFBVzvYR+2IYJAdIxise7huCPNnJ
kUGvQ0DMFxFj8aN9hdyGh8HeP03MW1F/E8RRfCCqvH2iaR3JQRpaBnrRhyuG5/7b
zIQbmkqF0UC+El54aFK05GpAcqvk1Qh0G4P2nqOwdePD6+yX6A5JF9C/1Eep8Rds
nmg36rBlcjzwQAhDJ53rS17PirlFNP/nIuApScSQPb0Un3E3R1AG3auq833KhyCu
vrN4wsiGUwdk//tCCdj4qZjgG/eT5kXoaVXnWRg53JMO8ewe96H7tb8AOEn3rycw
Q4IlS6MgCOgVXG3ePY/yPTFdHhAodkOk18vk2wH/Qy79f3vv1vglEwFGH8YzkbiA
h62VIrVg+JAthTArnAhLYz0zqBIxjHCENdS2WiYzZNniuLY3DDhZbkL1bRZk3Abz
m2OVeGmUtfXIRECU8MFIB9IHm2Qn09q37q1qbiViqJ1FFUm9O+I1ZA0uv0Kx6dzN
e+JpdyP3/8AtoJ87WaBs7544BlR/WgG4DmbP6KqF3UmUet+7imwD7M2L+/E0qnVR
t6Gw0SX2JhsI07vBfbCqMcY/X8D9l8tDi2VzsvYYvXFijp6MKgiXvTWYXWTEToce
TdTfY2YhpgYKo9D0M03xMPtoJnJGxYYqBQjvs+yatJ//ip2WgWhF/hExYFzYm88S
TUfn1/Oj/NbbrQXnFx2sCR9Yh6+9+mX4wzEYcgiidxytea54VtMmI8TmHef8uB9p
EFSfdh7TomaUdlktH2YlSAIw/z3O0t+OAodxuwcQVsEqjdNsiDVjZ4yNleohbRIO
8YNu++3dpYofCsTzAtT0SSB6FExCtHoa0D7YzzG8bvH+c4ctkWlu1Y/rKVyOUtqN
2QcOEv6luYDP+vuJgeW7unKfIpC0qbHEezvoxl6VbK8DVwGPtJ9IsHlO9VYzF4Z5
UcpQRyzv5vTFn3MSRRqgspUIIqqn1GxptZxd8Vrm/SCQJlCGY29RMkdYB3VMLViw
kjoEo2xfcYEZEVCBnlqmgXjnRNqyyuM5Q+QAsmEv7gAFdNYz6ic9VZaIbe/TDCo5
yakYIPYLJggmZb7I3KB7F3TCIkfvBcyjsl7bDFbW4yFfFg9if/TifTdY+yXil5GD
Cf8EKfYROYfHn/bU+Wo392zlX3mHnfT5dblxXfsmdzG1eKqbELh8fcHznprYzP4G
7beOuWRJHoh+ejzDmD3YJBJFQ1M7KaiZB+qZS6vIG32YzOBgkMmLwBrRP1iQx/Kg
Iyi/jERteKpewWIzA7zCRNihY/SfnEQCjI06FvSo6uZ8/qaYiOBzfK2/89l4NJuR
QAguZwir3Mqyztf2QN2Ol3VgTUokfS1GZHH3m1z5l1v3qv65A5B3jjvzTMOYMrb2
sWhBbR3DXtJgWBnmhFBrl02/2CKWJwaXynihkTPQ0Yc9t8Oh9BlDG4mmfedmUOMr
HNAnPelyFwhXmBFEyM90uGG2cbWFJzowEVCYMZi3LcAABNOwmZJdguZOXmKIHT7+
89/+AVS0A/4n3WU5nINCnSVIxa9qK1MXU/9GMiQITIuLaDYkRW1scQYDxBs0OwJJ
KgwDuRUbChlhcZgjn9rH0LVRpxyOWeKpGQcgBX3vf9AjH8I8JiHTeqn3cPSj9lbN
y4jMQTb3MHmAiZqUBvHAcXt+GRljjURr0P5BaHcF54Ux8uvAMRoGH17s4/3tErzm
VXLoAhbbi2P5mZRLnPz+Htl9V1xoGmNhCaOHLx1h47+eNlgtslbnP2lCZ418ne2C
h1MUGN+OwSzP+Wrr8fMO5+DzA0v9W8sf13mn4ivte1Ru4ry5Eia5iF8rLNUm6pn8
SXeFFobkjNjrpfykcV7WeikeCrcbVok4HrgeKU/MPwQfRwTeH75vB1MBqS5SThur
Lvt9OsWNx2MnncUwu7tsjNEtcE2fTgn50dut8DNHDrhygLfkvbD7IZQIyPmFnpOz
sq4xFzeu2T6RLCzTkoyR+iQIqikR4FraKljEDKiOJusO30M0sSSzyI8ktJOkpWll
rKTBM8x0Qpm1DVNakMElO1ox8duh09V72s1xNWC0r+Is5WxcBEH+f9nQeZ8rbP7x
ykFsdpd7qG4kFg0jiDUxt009lfiI97aOEuL3c+YGbyr6SIUD8OyxVJpbZVfzpfmj
UEF4NbDDnv58fcnQWogIRv5LK1jYS4OkbcAdLDyhL5Vib0W9hgPTQcKJciKNFGwb
ftgBO98cOYxdPEKflyFEg2QRh3oaPHahz7rYeWIz6wcYrGNEkxKH0rn2btFyj3qY
txOvMixMjZ9owqS4BLr8g0t/tHR6R0jr/OE/sn4EW8iduL3YWcIkjHu2ruPWsbPu
oD0tfYvlAlMwgbpo5xeEtMBntTm3wLsldHldgeaIV1b8fHLuUq1SCSuEj8Ws6qH6
y0jwn8q3G1KsnmUwi4NWWGT4L0LrxOJhqZwEDvQMh+62CBtjnM5PBcvIx+ph/5EK
9EWAel0ZOcvZYGzKMUKXbB3A3XeL7PwPYi8Du6KEz3vCk2L4YEkT4F6pjvhZm/Lt
Lp1dHBr7xb96ZRth5/gqrS6W2/sYJ7U9kIj1etDsulD7yDYjFyb9N5fvD311gcTw
Xq9+XDbju0dTi81bryJFz+Revm3ceDvgESgQgRkwq1V/Y/XFVBQYw2Yf8Q/C8aST
Wqrl+w+rZDiuS6EM6+x2Esql0Hyr5ga7Xe1upH2tT0OxyxkiF9Yor/knG9SRSGPl
NUtiHT602CTBOJ+EHobMFF82zcqJ7YWTvSypHP1tnCi1ejFbyjnANdoMt64MhVL7
lZJ/RZzMTbX3UvR3WmSNlaxb9Yb5kFVgkhd46a4y0nOB3DSIfr6CA5QzJjrlsizt
5lKSLO4eil/Ki8HQRBRYaiTz6ZNVP1O6mjBzyyTkk0ekilhuLIbo1BZHEhnbqMVu
HIX5y3Y6BcUas5mx+nhGdrZp9P5/GRypoohJzWWLP5kiwkzuhjY+1gBH/kBnLQQs
2rYFvXqZvfk69ThFB6zFTvwE7XPYWLO4qRLUVEXUhQLfkdmvAtIu+eK5lOXVtpC2
7fDABBcPTNZmHnrb5dtiOWmBDhMitDBDFkIhj3/AfSQkfUCQaAvukvY3D3Dj88kh
XFGQPZyEOnI0f1hWtRgsxUPwICGJQRMP38UUZHURWoGt/p3PBvl8icgQXc8NDXYc
AtC6bPGO2MkWg+CbQqF1DZuSuOd6B+TV+XxYcjD+NdgycGuZ3i23uGUlI9pUPmw5
ZAqHtXsUb0PloZfSKFINHXhWdBuilrZmyNsrYIfE9lTGRyJoWO6WBp8ttfATXpEZ
ghH+q4TJ8EZUI18RFU4a71iCtCjR3oQVuFAClChbXCY7GxfnLO9rT0oV0aiArvZO
vH8q5iapLIlVEXPbKn+PvShByCr6pRXPQ39VIo8Qriivdt4hVenuuhCuYLSiQqZK
iFKqaq7+FmfxyMLzG7/b1ulwTSA6IG5HQynPWLB71I/FVi4T9clATpTvtwPpFKAR
2mH56TedJ5R58yvgtRofZXFj94B0RJM6qtxCrGtghjhKw4yw7fTHS1A3G2JfQY2g
Lj0hdpdMOIObk3sk1Foaj+1NpL3QfPLulj7/qqFOMz3vvG22SJNl6TA1StJgZCHL
HHxKQwG+VweLmGy0jOFp0SFYJj2qMp4YYee0lFW+VPJ4stH09tc6/JyHR4IGx0AW
Vbtlwf0REGeHiS5g3aYW5RwEBOABv+o9Frr3laa50QVIrqu6PeIiHwzQy/kzeVDq
JGn4amJS+PBbfpiapa4NSK2S3Gx6QRnVeQlIuiFRWkHAFLgwJsTB6J3HnEMrINGw
c2xBk/HMPJjybYXklEuiBVjxdbfALe6Qw9MXFmHT3O8hLCLlmjQCZsTWm6wY1VZV
qLpzN71LNNVEE9mpNMruhnxnzfaOxj9u7WYjozbrbDoY8Gc/VTe4WiT1MYx2KaU7
D6LzD1zUBKCM9Q+o7W6G5K6/hmAg0nZL6RjwqPqbewDts0Ttag6q833zzHjxisku
kPtQYiwNE7E6B8iKpqEKzSlZfNELJLUQ5CUlJuunGumv/7LsbCtSkK7rSk2KNd/I
hB8R7SIxNqe2L8Bt+1jKzqYfi1gtjklZUAZznPMlHdA7IAUZXg+FdGr/hbphfRLq
1909hc0q0Na9lVK4vFY7iZfB4LFcfv9jL3WlHmd8VmEOyuaeHVwZXNGtksjoT2fX
fOk2Xv9rJI35CTzes5DG+VknRd6LIXgCymLcGmwb2FAV0rdMoc+3x6EDJEixlq4Q
HKVdn+ibqUBEkoDrVZi61+AQkTWRFKmdofXcHpiBSxW9nwN/CVwg0UNWuWL/ExzG
4R+NpMCl8X8CG7oXVJUKpcGtWSOyQ1vMHCcsqAuk3wDhzniq6HgchlpRWwxBMrha
dDArDZ+GoaopwHaO5KtXXRETHWlg3RsAzm8bYX5PezUhO2gsv24v4O+8VLdczXq/
TrcIApAP3wKOlSCQ5ViIqhh2MWuGOvTDyCO7m6T4xA9lQaaHL0bLXuM+WLkqvRXh
myGntJW6O/WVl56ZdzcHfzZCDRu3WPDZfWtysDFw0tulu0ic+q7XyjqUdlc7x/Ac
WQ+lH/d78Jo/MWQmEHU8D3UpWFMZZPdIH0MWYGvFr1YH+12QnLWLQWdQJVuw+L+f
EHbArMaXiEZevs44A3u9G65e9X7yyg/kBg4SoR9FLcvn64iB28PVqshmOQMh71q7
b+VPqM7Ud5yzYBpmN+0rEOf2/fzbSN5y7Z2+N3DJJvZOkUVbY4sw0kwySP7rNXEM
mwwPOBVp6PeZ0KSsz+0uQQdm2lMXEDcOOPOvzxTjihRbgokT9Gd0GTAgLnDvUzoJ
i6dj0TclrIe7hhpLtbLo3c7q7Es2IYf7BfWVvrpGvaefs3toksvz8K1rRj+4HdOT
4j71Hd8J0Yob8sA+229dOXoUdXlqv09I6EZtWBAaSdzVapQP84ojGEXc1/mfxnQL
naZQ2VNpn8juFZ5PV4OFq90O8xyi5H92wZOKLYdfo08uu7tYEWC/ECWm2/3roUfB
nbh9uQJJSB54yZVfZi0OaC3ymuhUrvYjHdACR6MCHOU1lr28WoZoerkNUFx98ilJ
z63CA281mNfCvbUVsdErLH/NPzLW0LSUK1ggTXJuMDb1Sl7AC4gBgQs7QUpinQe4
uVuxFv6x+L/2vhWcgfMgKJig/lu3WqdgtVnblNyuS+U8HvqUXC3MajqAXziU89LT
Wjjd+v4/but32+TGHHWW/G93/MX2SuhR/ZVzk+SQbGcCW9MgrOvj0IgiGO1bb+jF
pDtLYLKSCZg/JLfkEsqEx9UrdS8+2g4VGK2LF4OGBlv+gkKsAsbhILSduqb/Lvdt
VPp8Hawx78EQnSafTgBcR8ra1vHNdZuzTuBWZjUWptoXHvUG3OpLrYn4EoEfHmk+
Wv17KhhP3wfdpzFnl4Mye81sRv+aCyt9pu3uqyw5MkRLi11pmcGlIFwCUBGuR2kY
+vvXxnbNMUsdR8Md+YcimBQqeaUpDQsf5h8kpc/W5ZTudwB/4kEgWA7UKNTyHqfg
/XjNg0Wv1hT1MyQSXxjVX08h2YKQ+68zjsT8dPEaSKsOIt54n6PbTx92gy9/i5Lo
Ftc0bZXb2AkTNyFDpT3TqpBWZYsffk9B/sIWvP/Dj63NT5CCtCxpkpsIXSJiPs4z
+2Fsd9Dcz67Q6J+Z2fZlnKlfW9N9/H2e6HSUdOhb7z2Aa4RUkxq9SiaEM52UAQaK
p9Fgd5y8oQOk/kf7f39PzGjnkd/bsunTVah8yo2LGyXT5Bb81mDYSCSlYJ18JfP7
e28O5Dtm5urhliRjWwWNhSliK7MDOVAZ2GwMpLhPf/B8SpKTGPY0OwlxpZw4Z2OT
p5LMiQa2ivWbJr5RErJRwAFHnNQ+wgEmpWiNbyuGC0NQtDlTBmR0szA47rfusQHn
YMdMH59SEO4bQZC+sPrR98fHTVeqpKNsxC21WWr82IRZQFO8+/UYnRKe49jJjajN
eLuCg5rK0+tgZDX9jlr5+kOmSfE3JSdMCtttC9audQwDd7KY7rdsptaCsn60Izb5
sbcb/6n8XW1SJ+fCHqcx9FZjWvyAN6E3TNorPsEktrsbN1n57n8KraqPDvW1Z/D1
PfGfsoXgleU6mtkWZK8IftvD37PuKBwbm+zRkX48x2XJ8Mju6S9k5Fuqw4/E6Vt3
Xrgd4JyRmL8WA08Ic1R0H85MZ6es/4GTC4F4JVcQbdv6l2Ow/JmVNjW+RT9Qistr
Wjx6r6EYesbgim8Lx2k3YidfMzYNJKJ1gipe6qyTFtYGUE0wZIa0eGb3gUB3BGyQ
dwlBKh1/+OaZb/CB+AUmMj2VIvSQFRCIw+It9pyuwBjn7v6UnNhLmosMBhqj/fbY
418wCTZ/s0bIJM64nNTVNNzEXnlObxiAk4LymMnlfiaxzvvzITuF34eefCMl/YMT
EIwhm7ZQ0xroZQ7JiMHL1nICj3UoDK76N1iyJFDtCfiakWdU8rI3OFvEw/8SOaMu
cN3S4BELVtUPJR/M2BfsRnV+JUOwM1qvEWqundJnOZuTUT/SWdYPNEedIfg3Mpnu
Ao0DN+2r1e3KDZjeuQd8w7BxCO2XoDxIyytBqouTb2tXPd0XO1gaac1rkKqdQJEM
4IKbLS0PgX6EKTV3q8ylT2Y3VXqbqScUbh/pRIbiCRwjCSA2ExAlFnv6+DyFlDpt
gGuqScZxhaV8C/IUCTScbmtG7aMoL9VvFQouWRRlD3yf+SghlwII4FnZg1T8d4ic
7SYO2pKZ5U9Dga5EBmfzGz4kls/XL7eILYDvDKJ2wZ/LnJJfRhBJKG8b/UBAjGlY
embZOLYa4BudHyw51sQcQxZKwjx4arFb6GnfyRSF+9Znm2VkDuFUZpIEdgBvf6t2
w4APwRUbPgmrx/uv9PaAb3oPLH1XB6iJiOjwkclCfWKgg2w6KgrE/Ai6AQNftZtq
vXQMrHM8RF3c3YhJfHf48laCt5X15bl3cvK7hABTAJQ9v7wcvDBT6k0XxuoX/nlD
itz1n5DjYul4iNyqyCk600bnXYyxGiCnta8GNxagi9MSVLybVRCgOyS5DRFhSYoe
pVSYEgw+ijxwOkNeQssSY9LStGbX+L582yUY4rt1iLKqIkcB3g18Wv7lCVYb+ECR
6vsv4uVFbpSxgxev7TLuhQ5t7SG93ISytJiEISto6ZXHZEHlwr1pMxGk3asQUu/y
ts48uA2kQsJwqJFoaihWBBS704054wWFL8FaFUE+TYQG5m2nr3jswmjGnqQyR9KK
S5x/ZkBxqAZG6WVXWoNIzi/I9BwbZ46jhM37+PrfyfRbYYIdY6+2kruw3ohmE/Zj
yXcYOTRCji+3/m4EMfd1/6UILs28xC1ZFpJnHbRH62bTNe/3JBGUm0TBACsSXMQw
D6/ogQNF1/rliGw3wd7bZdABSx+bJb2fxJROtACJFsUdUTbjyIdMnlBi67peEkMA
JFCjXH8Jqmv5SuNvYgZPqY9IWatSVWqGCx1HwZZYV3HJaViywU0BaSS+uPWre/2F
LneAcTqTILc+59MYvBQMZzJCiPbR3P0C4KG6yjmWjL/oy2T3Kp/Zw5vjq5ik8VA6
Aiblm9Iu94uDrN3VgDYGYVCDxmD3VVwpHqWGhzomHgiJ1UabHHSQwSiyD5mrDTAu
+3GhVObkItl08kO3OWd138uJVHX7R7NYw1F/eI6HT9nElHd91fdjBTbooPa0enKT
ja3yAKpovJX1BTR/p7LLc9FMGooB96Rsa05H1QWqxSBMbHrM/0rwl38BmKV2qUZT
gZ5ND6K7YbmnqlVwRa3OXxk/tJ05T1jsd6rnU+VCIV269RXYpd10Vu0bb+fAwCO6
4V7arTABMD/7rudRPWZW1Cc3Sh5yHecwtBec9z/o2K0ft/MOFKmfpd+rLZC+uDRa
9VN2zqPFcKamQky5oP37kwy6bD1Fg/Xl2v2G7ZFyP7jWo9eUL2SWOydu0YbZVPNB
1TBb5aGL6UuEckuKecH2Of3jRoULA98SoLzRsBVUB9jqBEh6Se5sz8tPD6RVzSvU
e3PM5e5AfTN+S9XOZOCGEOY9qWoVuzTtgBpfwKYMRhV/dYsUCsVnk9fx2p83JeXf
wdcSoe5MPzXxdtRDFEHZP5OQiyyrc8y6zTu/CBabfa+KurUSdoAvfhfDuSOijGNe
GsVdYu+lDhuP8h/oAXrK6La6epLB5vSPb3N47SMkoNmE4SeEBi/8NA89Ae7QdK6b
uBpYGJdAbBs3liZpM+eVhdkpZdV/qgGZOT8e/AsJqAroF/czO2mtu7vHRrGEMduA
0bDXXbbt4crNYZ3eGSBQQ0c4XtdEhNo18/AIns65vC0+TuuJXDnoy+YhOjXTfPLS
JHgO9CC9cET4/4Fd/fThTHM4+kSSCQFYIYi1zggFf+SXT0X61QWjzfHb6QWAhhMH
2i8/vcT7mfrFVX3YAXpjqtIQFBALc/pKOwrIyw0SOI6nn1stCaYNyO1TpcF3TtTb
RBIaq7qFEk16bBTV7WFcrgNA5y9ym6JW2d1XfA/9o9Nsx0XVYVuMTA9azK7gFQKz
53PFQobQ6GOycDB0lgcy2TZvh8qVHbEZ+JQThKA5JwzUr85UDFNhk3910WeIG2xv
3/1O+y7YeISszYGfYZEBcDOQbEpz9ZQJ6Iw8infXMh49tTaIDky0LGDtwEBrrR7X
GtocO4cz6qGRAbLd7YNYKvl75DjjzSIcCIFP+5g4mx7dv/jv3BoAqRhN2NYHXCXH
K3LhDpW3c+fWGxSsmdSpoVDRAjLJzr1WefPA/vMoqFBedU0B9Wc7DCif+Sg/kfD7
op3o5z9LpP5z5OHApWt7WMQjdMejSt6cNc+0tTCsGiJ7ZUdRbynPF9BFQTl4zO8P
6lN3GebnMAL3dJtBamRaZWWEujLdrMH8q0NmzeDMz8sA7vh+po22JCYUHFWZx9b3
aPRN81pwTJBKz7ONdCgczRruTg7ILTkPZB0kcZpNdyhjbah6DtN2xe0YnWHWjLVw
p1XhZV/tzWSgjEOxXyk+74Br4toDB8cfrAgIBLdQr5wVNRlHF83ispYO6ALZV2ep
ugBU2Frla5DBMpktTt/hQPpMhZvGF2fq5dSvS4YiHQ68lmrlSlVGEPfmi/rBYHhJ
sxDyNED4ST5Uhzl2WVViW+qUqHMkZ86l0AOLZbAnFosD7tqcWfBc/QAH+npjWlLO
88LUI//iCDGhWyqHs9XllPBPVsyrtNZiEyb3dep9N6MCbsLKPArj5PxWXt6uJv09
dI7n5mqXcS4xfihsVn06++ytWvG+GUOYMeTpKz6C6S3eJxxh4i8qss9cjfypt5Jk
ZhBVosLBLCWibS1Oa0tsqXlfUqIatP/np9Zz636SUGwZtyDd34p74ZPfBSN72NSr
xmIneVWQfnkedQuXZwbHF0rh1mnVk9HbEg+u38NLhsNrHwBughzx3ltls1n+7SG8
prk6g+vQZm4E/BhZgHS0St45d5YPTgAyjMczdCJ7E1PpYlt8efcNEYHOfJKx3TTZ
Lvj7ihnJjT+NZSxXAXiQWzC4om9SFr99mD0Jt5Or+r+ovcB5DjwYEbL8OOh0uvRu
MOpLeIqYuLQD6D9daTpFxVl8q8BS5dEmPwspZMfApirjQr99hCK5m4Fq68P5lfdB
AoMb6AI4QiiMOdAKMyDOiePQh+nh8B1bFvYr8iHwubvaGGa4RJol9Y0JT5SQNT3a
qva9gXb4rvuKV9F+NADyDeCY68CdpFJkcs6MXLm3T7xNitv0lK9Ran1H1TR6Ecw7
r01sTkKb77/+h/GwiXm9cbfj96CzOYoFLw2tVVZuPyqESUN5wJcUMyILvLVpHZ2V
cmPhGPxm0pDticAXZ0/q6RkGMVhYRrVBXSpln5AGJOMhIbqvS3agA4xkS3CGyP5c
crBNvexpV/4YRGd/Gj4rQQFBZhhYoKbXaic3ippZTF9ln1QuNNSEzBdgSGrDUPkM
kWinkXA5Ohgp1+J2J53lTKpEU3A0cgFYqPBnMXtaCis9rA9O733P9p/hDiYTEI20
UBPJILHPQeIYsc0dDTN1C0EIk2019gEwsXQkCWLLL+wVw0zh2EQXwCusLWKxkCQL
PR3knIakwktbl44VoICt7IlxkS59C1Q6pPj+adg5h+PBtC8PkMoVE+Nanb3KGRk/
h0d4JkXgB/ZaSVLV7CQB0ZGLu7x59/OJ/p2gN3+N58psRlskjfEr5dalHaaFKR2c
dR+Uj7QqF8V7/DKNsAe3MkBcPl9EUhLJTNGwHlPbuMctGUrL44uquBuV8arsCGP9
FFrTZPd7tYuQvxgztqquaM3Hz4AbDwbeAm2B3uUIXDSgewr7Mw+2CqBK4A2FD3SI
KcgpzOWE80JlnSQH8n5V2o+9RfueBs6Ln5yAD0pGEJZznb+3/CWYysBYIw2raIxh
csra+g+zKnd0ZJtv18CNw5lqH+b0JiiX3zV1ulEvbTuSJG1umw+vkB0pH2VXhRBh
F8kBkZKNql5KYDIkwimVWWhPh9SDX7hdLaOSu+Hhxs9wyba+/lx+SfAMeXUkZXgs
tbRf/nGlYTb93npCiTAK7MwP9tuyq8Fe5PSLK9x/fhN2QHtAFHc8WrG3stqenZnK
d/BfoRxydnqAERHFl8rIs80pfMOuvmUTwaz6SYbo/IygYgfb38ngorRhFeDsX5aP
om1HIPl2DA7Kn+H2liQoprhaWXNWTEW+B6lE0zp3vnkzHm1m/yjIVSBWaj26F3w+
zHikxTDvI5bxd1HBXUk/eWI0bD93HUE+ueQK+uqvyyy0B8uNhY7fm3Sdd39XyVVY
uwswdWTeTjUmGmazbjXLf1Cboiu8g2DqFjoCMaCYlkiEBkeqZBg8kxlFIPwFp2Xp
axj7rpCspehoU/DhFt75pc15kXvtK5vFhOO9NL11vJCSfbf2qAiu83jQJaEg1sEE
cQ2J55VhRtb+7Le5n6vOHTHPGS+GWNyGLI9RmSJJgqiVWTlOgL/hVRhdfpGcWqMc
a8BCcb/RG5p+PdZKZfAGrH0Y9wNa/mwcSFbiUHQ2oJ15o4d4Jpr1wVkWpmWCmOwN
MQP44WQQhrmoxZwegXGer+EnBlNFgPJfhDBUXPHy88F8TgY3HK2WESUp/z4T4boZ
Y+qIpoldkRy7wMGHwcjbzxVFnTmKeTYvQIQoCfpoNWzwrHbAFBqNsmR4ze3pAspx
7DwHV8+vdYk2VCP0wil2SwUQ96Xym0hw79e8I9qajXggpP/Nm0aHEZn4JS3j4InH
LnVI3wOhSLeXnwIN/CuS9BK7AfRV/fNYCbquBORdgDLGXv8A+qsUkzUUdCQwaqf7
nBOuCIWapxAVWlvjDO/RR+wGel/iYLKiKayVw46LkQKr8fOP3dKzZee4bZ6cbCjy
4QqEvrPfPckwy90Qq/dcEew7MxtYVJszR1ocoY2KyViXsdtRaUlJVUu7f0WERnbZ
pkmrRxGdY+ZqNSok1NDoQh4RZDsMJqHoRXS4uG1Yz4IASLfRCphvJ2dM/To2b/KJ
t4qky3r9u1oZfv9G3N9LHM+LgDYcYhccKI4javcb1DzTRg5jDmbATDFZpw52QiJ3
kFeEnZH+/3zGcDjciFGxQWSIfFjTpaQDYcUcEaAACeYvIv00fER/ygK/yjyhhtqz
b/DD8Xslvf1jr7Whzst9vlFoMgoHtnEtzlxnCP+scNCpSswUxOubqotZAAKJ3tTU
ryJSul6dyNBQUwzGZmtiaiJMmTj/go3jVHdoAUK8Ey2le/Rnmk7QsGbGXUhXwrb9
lpN/VrBBQYqedNNVuf2CIi2qkPQJibVoJy9MMOLnErlD3TsDIfD3l4wIUMHnUZBH
XDnECO6Bs0m9aMw9ck/IvNGQ0/3N0QhQwrrkoFJF+EyIYFUqf174B0DjN9ISm9vw
7QkLhXZj1zuOz38DmYKLSO4CYPVXc9uXdfRFo+h9kl4Mw3FlnSxqcA86PVnc1NSM
voiRCsi2oIwq1srCjgtgaAR4VB/I1OaAkgbRH40Md7oz9SQsjgoCnbvLviOYyDmb
VNYtraaRQ++8HoMtISdcj32Xh4Kwe/t9IUAIrX90i7ela9XQo3coBHidOekwANoh
/vpIEPe3ePB43GF1WflelBL7ymadGfGdiWM+2bA//Tlk/rXv38eIJCdytUlC4mz7
otfytWa71m9j1pYG5H3ftMwFaoUcSEmzPoFppbHpXAJP+rQsDrl4+nVNcMWbf1Ys
BdL9zsYLfKNtKpQAH9oaSTCEOLzysjsxB5CsneLwNzT3/lIvoFrapg3d0/nxoS0d
5O9yZjlUNexxrSLHs1Y/YO3iUdh9R14Y8RNBl/FEH3/RQoPidjtoKeoBVPqh7RXE
8qheImKprwNMs0jUes6588AF0k5ciLiDubtGPyyFv9WH/vOuNAIaZZFlgWjjrySl
TwW8cfPbShi+6jhInDAHRmCVda9lFPrt5Jwdn0r+EgbUg8MHCb2qYVd9dDjmrgzi
feTMNNH0O9WWZbm//Y0zElbKNujaGy3lA+hK8LVFA2mAshc1YgC/VUsV+0ZnVndR
McCk6wK+qD+7rjG1s/OAcRhd/VKfYPanlzAhHr+lIvK6HYEMmG89ZCmoWsRJ6Y+N
FTcyARbLEr0YYZgYxlSOToptuIxkrDQrY6WHbujOfpRofoEtozctmy1RqWMpVs6E
EIoal69CcjLDx7/Q3gPXCHHFAb6hGW/SL3rmhzzN8zJjef3zJOn2vfVI5So2HpOe
vyv7+XM6vHh1Hj3zC4O+7YsTd1vXS33WF/DUuJc4vNQ9y0vzyO1O7bA/KFQUktus
xtvLMUIdr62LJjnHu3mKUlRTLg2l9NguO1hXYZov0kjQqGVcEb/eao8bnPQ/3sf1
M2Gc92HvxkIoCDhQUtiW7SdqNMe+kZdQ0DySTxqdHv2c+B3M7ll5QXD/nlFBGToI
wT3wn9Lm/j1WfKLD9WBdDEwos2E7SlBGb3e8qAHM/4x+7O7IZi09hcymWU14MMKS
DqGbo+kt/cWjmOrYjnEu5IyW6fjkC7+bQd6N57UWce6i3U3y/pFRqG8XtvjtB0cf
zYGp5qqvFokacG/FjTR4NYiK5mW9l+QgpCCJCmogd+Qz4ziLZvmTH2D3u0OJX44/
oPOC3O9qWHm2mfLLnzur1Gscd9TgmuIPamGqKZTncRimh6HfAmclF6xTK2uThbRG
WfGbz6FHldJFpfUXL7orQBtrhT43mHHmuwY3fjobqy3j6rk7nqNzxp+gnR2R/Csi
f+NfK4d0/qW24CQ5YZIl6dSu32JEI4RAErHiBPkOSGNfmyzqTO9tA8dFz2jOGBAr
503QsszchTQAThvY4JnX37qkuVU0I5jqyTqavWDTL5ZRQv8pJ+LF8+s5w7KOXse8
LAzfVXQ0g+sAnSwK7TJ9ZphnRY03hZUuw3/huN9Ex/R/xzbW5vo125QkLJ7Sd0PG
rpLaALxBucM/zDcH1G5WQ423dM2PWFaDFDlX5hWvR48mCpI8604LoJkcRmhEUvtf
4lF0JF0Ry0LnnDh+Bm3bDq5kvF1WZN5EFGyqAgSxuqHKFf6v+fpUKFXyL2k5hq8A
1UpX6bOHPlR27YbHVXJ8ai6UT6z4hZ6nT4suCT4EJ7vS5Y+NvicLViyba0dEuWPV
NrBntXXDCTlzGm+j2Fmlg9zIh/kDRh4hJE0eHfOAPaoo6kxu3QjttcUjEpZbta3/
U03Se4ZXQIU0MADqq2LIOH+z/r7YJUkqtaR6AyJx5FPt3hO8CTqXcg+1BYfZTJHG
ILJWi6V1JLq3oNdU9pOgZsBCnnpX+KlvES2t9liKbMCO+CdQuAP1FTnRGiNsGI/p
17TjZbeLX85FxEoTAfPqd/IrR5vJPCE+SHxCoC9lyzUUhazK+o8qWkcAdW6GSz5U
sZwus3Fz6VX3RMqxJZB9JzFERVy9I4oOVyUL/4cbD4CnvVLBlXttIJfXG1E/Jdgp
VeFk36g01rEM8i+zldRGDdEi2OjTgxhglojMQkBJHXIWHlRiO+C39aR5+dc1NWy2
DsmD9egMjkyNzmosEMfXD1q1TctnSTQ3FN7MHS2rrJPtG4WWz0Ikrqjo8qQg4C84
fr77FfSee0zTMpgq65o/vtsX5VBwzCeFN1OrjAwNP6h2vT0ZW51LXCC468RKvqHb
5HRzrVp4qTlyGeGan9FyrdMJPiAN2TfLIVXJAECudmFSmMXHMl5JYwjy8iOfRrTk
KXYetEW+DiOHqyVU8U7F6zdcr6v6fN+NQCbTTolEjERpOZo1K685nlJ0rv5s7fdU
8iUKwZC06jOwM1itlsoVnLTfgk+xO/9YaxuLcvDdxgV5k81NETeaX+RdX83wGPmA
mEbMY+btS6Sbe4b3KFfj32fPWF1khmyk31u6hATctMmY7cr8Hih03Cv6ACOtu3i/
UX4X8UcClk/BL3jesRpbUOzEgV1/i/tWyHEZf0Ggvf1/9jK6CmmnW6nBJLmorks6
tqy529EoPljmfkqMiyMfAB6DWhzh6o0zjnF5Z1eNBGo+r4tpFR8z9sayVFPd35ya
PbePw8/Awv9i4ajemRcCtTv+VqIRyn2XohLMwzgzG/UsDQlrqzEm6vkw4x+vmXRz
7pn+l8fqCc5dX/ckpy2ayeEpRQPuHeHkO3PG3in1ztgNLwGXQvvuINyT9neL1w9V
NgYOeRPuBYziD7XtZiad6+hmgipi09nrwz0J/qjJ7RQ9rFUKtdXPwff66Hv6xob+
OlUg0cFjhFSo2SsO9++NSehPZo2YwrPFmL+7tZI8IhlrUs/QSdCZOKCr+VKMriJ2
E3ONN/BuRQRiE/LfVUJ68YkbqAIZ8FXhXZaxV0npLdbSq8X7VK1T6+XmyKPgxCiu
dkRSpVyvMzfZ1+H3OiNVRJZHHHqHsl0sqqbQt0vv8YMxz1fl3Byj378LzoIqPPrD
iARF3sn4HU+NvSP6icVFhetgBVzx4kdcMGWqwVkcJSP85g/L/285KaYyzgnOIi+7
7vEDJmd8vA7t/6Tiude/Km+MPOpRKOsdRDP/ewMAaLRLdH+PSSe4+OIutFU7zYwb
OMUOPeIKcuL823kdg2CfSlzd/0z6iHFcgetCgFPcGT57dyk8Ja3ritKWAhKMoLpm
6k0n3+7OJSVx8UrvkG8ktAUkXF7oVLTXC0CGozL4Q8tp1zG8westFr6eMzez8/9J
GgriIjyuB/UsuNW0RSuyJsVfMpn3i9ObSZz5PkOv13JsgElf27D2A2mEoVAp/RH7
EaDM6PRO54JejO2KBf1OIr305mJkdkXt9SHWvNM/2dthmtY2kIi8szr0SVllpViO
C5McXCPr+KCxoeD/g4J/DZ4hr5Qm04tXcD7Bwv0r7sK8uAbQEkEjV5OVWJCNVTO9
ge1dwL1iJgSDG9uG2JzNfgXLSUTqBr7VI4ZLzAunv6/u+bKlx26jVoNff+mZxpT+
IwVh6OY3x2VsYlnAdVHfoW8PTdPAAfH217DIRs8XxDqz+22zzBh8Pju+jqoqznx+
xBTLmxAtjVbwR16uNdQ5h2hiiLj+X17juVO3klj7G+/2rjpmnLKP9NMHBCzPEz5+
occc/inKzF+s2ym5SG1GD+h0iPCcgLoZ9ST0Ue5N44F3/Kl4pWH/0DlPWNmMLe2e
OyDo/kiEZ5j7/1NUmbf5epESab4zB6j982JWgkw9RcjPNhldmza7d914pDGRomzF
em+yaSKCEEJXQiLcZBexflKgK5wtzhtDeLBJjlPmMCsXPGS5juREMnEpfhOmGAXe
pz7DAZzD0PVIQLTPzrrlvYDUwyjBagxH+PUTNmYmBOm8RNsMVeUX4wR+bUBSNb3S
GfU7RIxnP/BlAsqYgMUmd5rj1OMx9sEaGlppBlMS15AFJEZujuKpuy7RnSmsVACW
YnM+FaEt9D1oJAjwKLOwRB0fHGGoo82Z1CsIFj851NUsh/kr9hXMslMqORxXWfNd
T2u/PAfdQAKaWsWZut/bpDTaJpqXl5r7PWWuYYGyWI0HBGBlRKkwVCdzKhhJsqTK
4IT6KqCiZlsyC/BR7aJh6+qt/qKWIs2mady2bLevY2p+TO2lhIqb9E6oBvKwm/h8
gWyJLwT0Ymhkpv0t9ZkV6zGdb1MlRMcEwMJ1jv10354qw5NgXUfT/TzJyz4t2YHp
Umj0aOwx0Yjj2k8WEVAnJDkyF9o1bZ8N67+fcjhXSMBUXiyL2KPixHeT48/vkojK
2UZjTkPwIzFPLylC1wOfy3+7xS3kiW1QsG58AbsQlSyG7SwDectEogBXWfhvma/p
prYci5rz+rY56wVDxpTgwL8Koc3hutBWUIqIfsCmIBY7qEji0H5IZLRhztLP5H7y
c/ymEUv2ido3GGRUuPLXZWxy90Fm19lWq6XlMp3gcV7XRiabh0n+WdQ2wSKt4lF1
oPzT+yjwEMomfc1anorLzPVNIk8JdXGRDDJttwPuzLhQtf8egw9RkXBUZMxoBHhk
AGvVNDEVcsL9BLdroDLNOF4N/LXm10uKuYgs9UPNiC70tao0yvcS2UVy6ZfBWtV8
HCjajBvvqwyc0GebiHB8VnMrnNK/3N31q+Pc4b1hkJaTAePJl2tXrmW0odDHIBMl
Aut5aMKW1Q18F9pFvc34PrttrvjgMrM7vC/PefNSyS8YewHP961f0ASy9ySRIdND
+dawd+pplHOJiMdcDz1YQoPHYPeEqoCtu833FhmVYijHlDpOWkn8amiYkVbGgkxC
y7R2WbJqgJ7yCiEAmG+nnyUZHD2xCJu99kiBfvDv3+zOuAQok9sX4cB/N55qfFsn
9miNzlCTaZ4bstWEZruDNt7UfYMmcUKa0t/0U6WUTHvA2dNyZBPnMohbX3JT2AsG
P9Xv3Uj0aebLWOgk2iLtwdYilzRA+v/rk7q0kq/+4LMzrMdjU5c9JTNSb28oEham
FQH5OBM3gSLGfL/taHlAuRvTVDyt1ekGTtnfUINTKV16oIsNnsw5vyT0QJGs2YTd
hk4rUQJ/50IGzwtkMcQenxAogZCmmN+00ffcSJ8+P4iRBD/a2BbPFTLKTZStq8ot
wxXXv3EjnkkEPOO7bA9dV+VwgsQxzBRt9rpMA9b1t/GdAAabNYofYpWdTc/zazW+
QcjV+G5DWFbbmJgcyn76fepWG8Yotc8tMNI/WV5ywQbA9ivG/LWVNvr2DSNdOfRc
hzTvVO8x8JwCTH42oAER9CGS5t18WnieLlnR5rXevFrHPiGsdJ7mOoSRNO+i57oe
vcYRItNoWAkVDcFLExmE3mhQEvDZ6aH7gHrwmFBYibnXSUXXlOto/mPfPzTCj5kV
BJhAH/bCfuvWcsmsEMdIpPhbIQWqOJ8dkLGk0UUoElgH+DNY4aKxYs3RPiChJX5t
02fZOWv22Si5QyTgsn1ZYwP9Gux0xB+nkDA6gMD1Mg+ghF0WxC0QXiCPy+iEpOn7
P70ep0NYsK1o84gN2d5TrITgMBBp8J9qrShr+qEq6YL6/AhDYithID+aP7PInMzS
k6onlE+/2zrvAhTa6Fu+DnvgneTR4FN1WuLmsNKAWVJNc1F2BcwwtZoblDH0Z6sR
TjejP1MJtmsTq7A7Cwp4L33ZIUwv/QpFj77mbbsGsuPzGZXu1h+AG8YXkesWG9P3
kwQ2fGnmn8LaDSPtP1ajuUDuyM2fnCIz9hU0GfWkESsTdsjSPAQJCyzxnkCVUbQl
YZvZJ1TtCYyk92OFd9eV3kgL1qDL16OttT5Jdu+FiFHjzrEtoUe94lfFwxxx4W8i
3OF1UE4FbyvE2h9o+ZKToz780nRnPdTSfsL/VEA+HZaqj4JvZKl8KrldhsfX4sdF
nJLmdjyJR8bJNvXEdXdplnDgVIwPoEUIod5acpW/N0P6WqPkDwMLEqXHULz7rf7Z
vZNpGmcFbSQipsq+2VxyleoWzy9wm173NR6yDM6WPFIQHnoOSzuZnPAasFO5OJRq
XPmTfo3hPQlHiGwMSt3ctuES6fVmpU43TJgr0/Krb5mwNnX6OkIkN26847gLGlbZ
ll4BwdWoIcgGvwLTvR+iLu6cCAsDVfBi2h+h9rMP4tRnkb/F/tpauyIxjBbYwysd
TcWLpMRfNlijOf6wObK2UQ17I0tVst8qGEMORSL1V3VloYzJ6SYlcsh9ctOn5lY/
FCYEGCprAnfIU4HGlYDmR2IOlydNNIfLHcnM5ZgIy8vyaJJIhlujXVTkOYcAwK5b
J506rUmUPELgxHB4ufv7lycHXJI4gAybZIE7W0nXx8PmFLdH/pAyAQ0WvlIURon4
8KeXtIn893QdjbpzHcx9H1IpyMOVriKfoMnb/bUKZNHV/lMmIrp1WNpiJjJiMkyq
IfCBz1jBkk/NLnKz3oAb8iBMtbkRrG5MtEs/A9fWhJzCF1nQQbE+dF8uWbGLUbiJ
gJ313SzEZgQJvTPn0+q588DIotduPVZutOMdEoA4UIUIkPC9rdj+H8vRt7znbAhZ
TQzmVHosJMWc3hkItPNr4J2DWfDomfl1GjpIJGooS5b0K7ec7zmQqR/1Omhwc+Jv
PkchnPZM7EqKUYs2KaW4VrQwnndwwRW9kwDTSIU+zFXmilmy9gN2LM2hbfGOsu35
yT33UFv+CA4050Pdx/4ilYI3f+v8WLcYxFvFxayHkJnL7BPK++3AxdZ7+KW/H/4n
HeXjSrMERXMVMy5TKWbAnGDOHJGCKLLnIsMbdTMAu/N193dcEiw73mulIHROTRTI
s1RF6h4bCc+EVeSCui//D65h72uvF2jLBU3QinFEtoPgNI1R6xIRd65vmrv5Hwom
i1MSu9Dji3AVyZ8Wez6rJa2j1cmhSyI5bLwUM4WXNm0IrJ1slclbcPjRO5Rcv4mh
9gL3ZbFOmDQ4q11q40KJXoel+Yt/Az5f5uFEXKJxg1pFgC4mhtMZGaxnPufh33LW
Ux+c7tUuJoUB6OWM0s6o+v0mDAcQsYOkiszeKCaZQPmJ2v+wAlZuCrfMZmEHU1k7
D2x7/SuapqxhaJZCQapi5ISdeXK9SbQX3nRjFQmrcj2HtCmD38F/c47YO/xkTHdj
fzbkxH1VTxYY21hFDdhhEOWfDBSCLpH9PAfE1Wtkz3E7ulYK3j4Egv1jc6YX7U9r
vCYDjFoWJzDUeqCStk65ClryYYqYuxZQunVsgWfI6U9IYLmMu+8zw+gS8wnRCMPk
w9lAu/YV7xzMHK9Y27zK+ZYXHLbD8W/LGWErVfO4Oa14KtKHSqkmmAFA+vW9U2FR
W47DKmTzNFnEQmhDQfRfZWOpyIQZOUt2pBs9CDT37zCZ3rMSn+7vBxvoLDyqlit0
6e6Y9StOlrPsoYtIWtEJuz28lW1Kc/5/Bq5QzHp46LvKMBFUmo67Z5rXYTlrbq9c
+k/SBIf2u11clzePZAo7aumYGmVp7AuR179uGiRRuyGbLxf6Pyvnl4U5v72mLpLr
ig6GgC1w8imtkd2ePKckfNbG8Ww4qLo5ynvuaF+a/A5/X7t6KLfd1EOU+k9a3EQi
/Z87O6av6ITi/a2yhZ3ZxpoGEgRw7r2HVVApKN9DfKwlaPsfKZF1gtoB+SUBf8/S
bVREnfJHMYDNjyEBzDitOtCEUuvc7RLPWxqeI8Hg42CrUeGJ3mbJCPxUbFD8f9qd
wvivrU5jjCizOKlGvsXqZfxn5ZidkcNP/M9VdOLVT632pUQU+s4vcOCfgA0r/oDM
4hgESAU6lpiA3deofWHQDWtoD88lZdKNsgmIYFfCNUUP0dktcJmsGNAQBpl1nsLB
lk4w0CJg8G1MPr4BIZgDLXyBaAvnylOwiAbsHITJ16uxgtm98OHBSDylGZHKRm2V
iZtwIG0CGHlWbH7pmCIiLlrZs8cp7Dvv6QtgrqguG3eTgJjWWqYmSYz6R2Xd9PEx
WbKTzzefiuuc0vf2cGc2sVMlYI8Z+ATlBUKADZiGf6A02nfVL0KpcESivunwvN74
LhdiZepvkvHKiyVbwui8Z7QQw6hDkbIWBQL9BIMJfqxnivhmDykP0qIULcpc6F1a
JcrC1ey/1KsiUt9XLFLw4rIPtgYaNe98qHhSxd5nutD3TC+uitQcl/ZAkbchVTh/
PCdd9tsOBrq9sHDp4ekhSaImXSfoseH/+/cGIIGqPuqMiQQ/kTjw4aulfpm57xjN
zhHE7/ArxGWC4PnieMhsqt52bjr3JsHrtDy2wf/hHPTjMMRk21997XxzB0nPCW/6
j50DG7FRAa10pBNTJNBEdxfJ6JBShpP7bH9e9QR5PZWoHlQ6OpWgjQHaJh+VTbDA
FxLQp8MfVupPDpLn4HNK3QkvGVWogzsRBQPrpmTVvSNRr8bRsedpKCQYWUwt7gK7
9fCcvHD2VF/JFzA4Ol9CzcAmjLWs0MN6viSxMQavHN+VeRBtaYkCRNzQDkGHOC/t
FzwjVo/ALa2yqHv3YMxjN71J7xCr0s3cIaGIUddQephw657zPzBE+5fnEPGKBt7W
FUgMI+1TOSkZZ2d/GTHv2wpgScJ4HE6fymATFurIZhqS3IbXqlS/uQkebhFyomwF
eqUAG2NbhYo3fanq+fdxeD4N5FEVm/iwb8HUb5GxRh13/inX4uml9jcvFrDziQvo
uubBLk+wuSA6dH0QtE2iyaJbkfgFpgF5af1wWRrTPvD6Mqb6lomTbwF9tXsIJfKr
4K7Suh09VgiSUHSzsVsYe0W9phHRBFEWRXc/t8GKZ8I8XGvjpnG6tC5TewEB1Dax
P4HlUl/uu93kNig09COtf71cKeB3DaEFsVr7WBbV2unH74TB+lEj9tPwDcf0pmdN
OGQ5Ai9hmPtwfd6kvopNgoyOc0XuJXsqSrEFeQ6t1Yq5Rsaz36yXUlC62L3CtSK9
PPEXzb2SFA0Z8H498vxcimrzg1aeCqu6TXOWx8rcTHHoGu3uTMPWK6+3c6GvK8xY
X6kh91uX+zmGhohrnlmdROK89BgXUmmarEmBWuWcVLLu2J/r9rRfx3+MeCf9rkfC
LAkvYcrcy7iJCsz16fGC7KoX36w2cVQsVs/K9jJTIU0vZ2TTUoKbS8G0YgLquFDI
Zl0CUcWSuRAxBuhYzLMdfdiBHJmDB43LkRXUA59y7elHNcs7De+g+GqNwafz3JGc
9e61EJOpcMy5ks0PfrwwjN7YNrCi7KSpjSPU3ZXnlTrvORwU/AVihV0aW3qGazdi
qpNFtZ6bgueg64DgggEWOxugprRdyQpSZEj+Gs9Zo3h4A0KtS5AWIn/Zgu84G809
NyqtMm0XWxrnPc3Y+0mPMvjehyzGCP5QkhxwE1ShULv7gpc5NHtDiDXKxMd81w8r
2YKJuNzAJvI1491bSsn0y+nPyThv2jkDru1VqAkmwzCr0KzET9m8Od/y1+jth488
NEjnM0cejUBGbFD+ENswrkb/ma3onP0/8rSbaGWxdT1PIHtPjO3pK1SbdKacO0fH
aK12jM55wCNFCpTg+Fktkptcqoy+GRD8iXosK6FfRdsDVdmwYeqwKqYV6Y58E40G
ZOzPK03IJpf2wYIXwdfSDN3lODhgYPkoMAOd/sMx5OkissAy4Z8TGhmWQRgkiTBU
w7Oy3oqUI/DZRQ8bXNkl/hRTk9NvkzQ12pCBVm/0Fjml3RyCOgNqVdH228ickgkQ
k7iI2Dll7EMSbgAw3ZOr0Hc19YO21DkYkgpTcY/mc7tDmHHGCMbqGd0FKqhhvRmV
qkdwgtyu7Gd3A42hWuqYvHMRUeT9ljy7CYon6N/GsK1BZpWuxpuU6K4lnfr094Mf
nCLkGPOZ//ZC2QSA7ZvRfjrU7fI2C79lQB6JJelaaUaHqNkLDANvKIf5ITt3MeV3
kfhb2jeTvpwUIP1ZpBzoHqj5kflvItJ4ElLmDXz6yA22AqFjX8Ow22UIlW+p5X0e
3VxlMngEGxuXwT9IqKAbGV5WMINsljiCL3v0Rjm89hcP6zxjbcEchNgq1fv6WzPN
qZ8NuqWJBLwfg5C+SySUBIiFogovlp7KDZkN6GnhIkYpGIYXWfKozEeqkhIDsVNk
wJBMLvEOQzT7NPfTb5eOp2Ti9RdVwl2l5PeUfNVojD9LNe63JkcOhZh8668VbvPR
oOZcexqPzMC5TbDC6hyDCF6gZDaWHUzIkuPHOaaXGJdniSB5690HJZ8WzcvBsapj
8flOClZ0UREkEvy9Bn4UAlI8AtfHzBWv5bz1s0IYUq4makvPfmuUBXMS3VOW+MR5
EPslD7f8dvt0dlD1QuNKQ6M7T0IIkJVpkqxxkDq0Pi2Yl0excK5BOsutfjp7HLCX
9S6ULKTYmn4DdJfcPmFY/Ppz+2qtKZ32I0uGUpLIocNUMEw4ttFE3GRSXbydWS+3
w9bD8A5FK3PUjQx83vn6RJfaaOxBuq8QcFlwaQvdX9r85GpezMaHQUS8XCHJk5gY
TpXjh2i63BTvub3B840fcDET+Ue1SWnKB5PGBrWh33HzK0J8z83L7an4M09QBgcj
gKKLddmsS3Fh7m/7QmUFRlBI1Ic0Vy/NMaFH+f7FalzoO7COfxA2ZOOePmWXTjnz
YruVxEHaXMwpE5kfV1ILyaUYB/j2Oe+vklHHMQW+oLu+pVtvtrBy+WfX8VS/34sT
z2l2Sts4fjAFt68cEqRCWAoLCTN74l5Psk9wOZB01kLjkkKMfvCRaFA0JcxILc2N
lbYswGq1J5/+Xwdd6cgTw3PPAyX3oYcltWtyaPhDPBVNZiu/q0xM5lYfXele+Js6
aHgpeBtR7B1z2wT0B0FML3JvcCy+JcC96C3uxeirzSXTxNwwwJLgszOfF+ExRHbf
3hgX+bgfG/rYIfJoVdG4S1A/sijRwFEXYxzuKD1lQ+BHd73Eq+E5nJuY0MdB4FNt
BSr/pDULOEh37ZW7GBcKQbfRwQGBTLrklYsWT85po4wmZ+RWa6C4u0yf3bZrnY3r
TtgMBqtxoQP0uo9+ALjN+cb6RuSxmUAH/MGMrVQfuFN7lBo7EbkkhIF/vUFcILtr
ec0NifUy6ZZX1Z4IAgCam2Ml/6LQIwT01RyB+zHyECD+q1ihl4/0tkDzvYqGFhJr
MTB605K2x351lvAjDSSffseS7fUsTY5vESMdQTL6kGwOQaytIMx8s3K91sSGDZMk
pIRw7ubH9zIXm12EkqnwJrtFzumb0C1WRZJW2IYHefaBdOzeItr8bJfsMNDVmp3K
PbEAWHl/e99xVOIY9L9cvlWc5lFKRLmLELglxsstgAFixPKj3UMCEtZA6Fr3oOz8
AluRAi+s0tFWJdJkyS4FSAIwXPtM0M6D3woLZ+AhGkKdxbosKzafgNQ7yHDUHhbb
GJ8CNNSKWaaOSX1F0NAcor2Q+8pN5qSWvj+36PLs6w4WsZPjBoiFmrelAr8j2G37
iy0suj7EnLy04pRnK2DXCWcnEWP7XX6wDGziMx20WO+SV+9fciHIdAdwYKOKxNqO
kEncfUgQjEQ5RsxsuwaPuzYKxHnU06h3utu7olxhsxV4vmQBnuSqkFBFXlUSQFy6
3n1YzpKSh10lB7lzMir3nt0F/Qm7K/eN0uQOvriJlqYNfnTXLoZERIhCESwmEJA2
vRnuXt08+O9Y67Jltn3vK+PviL6y7367O0xoVihb3w4Mg6dUPU+1OGwDvGGmfg+i
f02FAxaz2pXa7qHe7SN/V1ORO4cgtGSQnGeHsyJXli/riEvdQH6QvFfMpKOtekAY
PhiawQe5Eu2cdMtEgofDIPJ4fScsenxJNsidLWCmZGHcGa/QiSCepj56U0JjE6hi
d+Lb4Wqt7chZXMJaJmSKaHxcuKQy7qQeRFR2igYac8y8io2EWRJQKc79ivSF+Jmo
fSoO9xOjmlzvz0Ps8mdRM2yFLWKOJrQkcd3VQ5cQobtIW63V29ziY5Dsy77N+4C+
hUT8nsuumihUHL2Yxo1ocaQ/MDcdjwcfNu3ywFusEpL10EFSMLpVUKrskTfXWksa
eV3mehoPbYsPrw6V428lZlmISv3ukVShTzYHlhlhtWLbH+5YOEYNmdl1EmlyYI0c
dFzSBifhbvAU8+YDaXw3ZeHDjOvOTB4aGAuW/zkOd3Dzskc/XbZEKW2LLETYJYa0
jdBdmtnKUsG0om+Xpq0/HQxIgqFRK1Ju5CdLcMLVVaNqjvkrVlEo3ccb9HRVnkjW
gSmwwW4iJBJr3/8tPEnB8g3jACRjOHISaeKcrpL3MK8sYZhr4IIfabfZD9xLbpZV
cs4hC8j20AQ5K0ihp97aWtdiW9bz+6Ht1W8tABeHFvI9tkLInjRU4Vr63UKdCK3W
chGnQibvKlK4YND8wyJyjJc+RdibagxhrfQABUERsBrFm48xv1K6QCETKpUngB88
3EjSesILodwWlHi1BvI6LJ+40Ysk98fIy9M+wD9bZgX11dsUE9wN2cL+Y59SgSwp
xxeYPDyKqfWMVsgAWzEL5DM1MNxzN1yYq3o/oT8oIfifuM1I5g8/N3Eap8yz10HL
lQpqbg9g6PiSCXwloO+o8fFiIgeuMXSUmstCJXbM2S3tMOedytHjIFaf9o7X6RA0
0qGv+VtPpC9pDNSqXv5LKjLp4Z+CjKPicnThwZpMpycKUCtSMW4F242bkwcGBSX+
6nFH+EnS+/vFg7V+JEjpg5yUHKThnCmz1BNsBDY3/P+NdGRWEVzfx4zzSegihQMm
oj0cfEsyhaWFXAp2eQwvGPQV+p4QL6lgpuf195p8deB9S7LJMyyUKD5XLc6Zkio9
XRMWfpeH57uZuuOpn5wFyHx6Xty2cqAaJcB7WdS3veBcEgL2iepgCGKoN97fxg2a
oIITW10RlIbpv/rT9MtEw55b0jnD6AWHMGluLHgfNc22nCnAOg7TvjHkRH2mflQa
kGZT9RJlFBnUfGMTigh74ftUkPJPlRsGWFrjwBKGSM3TAt6Z8W10dT8w6QWbkAuv
a1mzFfYFBLfafX7Oi2LGEpM8T2UzGSaWQ/a+RCm7iObu7of2wlc/AJ6wyVm8bqWH
8+gyMXTn2ZfcvgOj2xD+YaL1yDccADjf886R6ZHl402PBMGWkvFDurKo+W7N54K2
MT7tW+H9QVOxHMfkAX0qaHplRwSIul4jRrqu4p31Ns5MajsktNisR6FYJR6wbByc
yRp+J8FiodaKX1ccbpfTQKhEC2cFQFZO9EmLF4+CR2nFSUQsd4wS4tbhmt4KTFlX
Og1bLqNGL3nyG2NZbtzpMqasheIyQkJyQVZp241inVz9kWWq8vtlEud+T2y9JC/W
XqPk95nb4pfYzqU6sG1sNwuPlbSlrkk4KSzZQxW4qqsyUAiBFfZIW/opHVTDCufp
GD0m7X4C8jKLco2Wk3qOLF/iPyWk4HDDU//fw7w4CsC7VdXkZQp5e4iKHZi7ljRm
vxsy+/qXCIc1+QFrWKQOdWKZjGI+jBhkQarJjJmNZydnLNlkdiqBnupZDQmZeY4C
QOg3WxBV0vhz9WU4dQcl+wWicjkGPTHA3f/JhVxtsxrf0+r6tXSYft01zGp4zfaG
IsnvGt00fkXUITVsUvm2YfaxpL33KDAiGMp0HbzqT/MWHiy/2ycEJyILQHtr1I4h
1bZ5x3Dx4fKHNbCEf+OvZw0SiaLoFNDKlco1HFRm0S2D7Qm9IFJKNbx1jC13qEO/
+m5rZqsEVYySGW4/Eh7HIGSkXes0biGbJZOC2Lm6TxXEA0u1aBdrKrzCS9RTx0ML
pqRtRu1BjsTpznADrSUidCzwkbSeeloHIM4ylnSJMa6IfdR0SzWa32WB1rtQQ4CY
N0IxY6jgvICt0gTaQXDPiVxFMy/Yc/1XF3g49iiZAJuEdidbN6ynbAdBb7/SqQfD
wYi+j5YdWUfj+4hVgqlE4WtxzaBwZ49zE4nnPDQG+2KkSVInR3cDioJ/sZIYl2Fa
tit2sOX/m9aNTTwcdP7i+IKvJwho7Fi4tj0TKLZYOqpW47vZ1PVxISAYsHICH8aa
zMQw7M1pf+l2TFGScYGa7DEyfgEIaAzGkQRKJ2sWc/mXauvd6K/S3w8aiFSHgL89
BTH++lPSomLBU6xgfWjUK+N3l3TyQMLYI9NYMGb72TMY53UORUmaJKCl8K3fSGMk
/BBnG0PJdoBVSDExhgjct1I2MuRenABw+5fgpzHglBma4DorVQqo53USDtmNh6A4
200OcKCdoztlXXc+j6FtbajAOa+1+aMvu1F5i9imqdCS41p5j3Zn1eqbIrEQB1iI
nJMB6SGyck1NHxE1eRozH9rN+phgb2ROITPMpvAQe6PEWSd7MO5PRR/K/Nx7vL8v
kv+yhNvVrYAlA4za/MJaAQqdQIVCs2Hlb1ikOoqrqapSG5h5qkvoUhcPweDuWY1U
sT/sp+gHi23jb2BTmLSGiNjLs+FswRJMa0ehmBbQUqS+6qY4lngdAHsW2noIaEWf
e9tolRLtkjPoKgcuOSk4OyIMa8gMh5iicrAb10KIlGeGY+Hq+Ir0c4OGdxACNhfG
gbrss2MisjQStNys8xKfUKPQ/K1uk8Am0y0cUjlbx7qg7L9N5sABXAvWof7M2MB6
Te6liCXDIeINgXGsB2rn1GvAe61JOEIaN/EnN6jpOb8TzjysT5Bv6igP7qZPw6j8
1f5zSiw+Ikv2ieugD+bwOUdy/mhPemVLw7XDTdzc0Sf/2j+QFXyyc2LRAMtnazKr
reOMY3GmVs4AsxerIoGmOdqdLO629GyGDlom5StmJoF4E/jBCms+AtSJtIsj4neD
hhR5ECaJm9eqO+gekT9nneOW31XsLZHiAyx4SVcfIWctzPbMVRBfTsL2qCdcBqxl
008OCb8HdP2sr5HsFFgdEMxjropLzbJPwjwADxnzYeTr5TiiikFRTBaKjjMIAKD2
fMf8S40L/WpLVJtOdO9opAnKC0NsB+4a1XHGtePzGUYCb6wCilUxRAvTBPtQrXII
KYgvcWdcTkGHE5LAVetdGy7zvQxw10CerEgpeV1Op5sHsdabUHnceB3Z9PPrHJnZ
BbUzRNDcLz2B9ensYaGEoFnNDripIiBzz/qKbJ4eo9BrIkaWe/Pqc1lEpqpkzSSi
4HAFek6ZY7rz3LT8T/VQdbNIDYiJB54NwdJA1v9vrcMbN95tb0Indrczfpfsz7yY
hPr2r6ybrp0YHDxFwKd8Q2sGwo1pUJrG7NrioPYY1Bhj/18efhF554zVqMlr4D0+
RGZmBV8IRMDMP8UmFCrK5DJ5xBdkURwoRVVI7z+l2ODnDZLm66V6cAYV4KNNSCwY
fFy7qONCTJ4+25M88a2LXA//0wCCiDI82eBxCWgTDvVZFFYJMjb+NMoIg9kEtu75
u/25wUyueOnlPktO4MGXvFavjRHXLr+BOsio4SwnPn/uLWgXk645kucPV9bqs3kI
WrjJ5NGKb00LhJCFhwBDlasRrTJTJ+wa7zCPPO1NNr0peVzvuRhrh70pvnOeO5qt
Ea6LgL7lQQAAQZUreLsDkta7itlO8nEOW9Bi8Pr62L95togyKKGiRIPuZ1iHIrBy
JfOb7BeyYeJUUl28438uzZssvIqkv35Qxmv1C7YZTDOhZLv/fg77ddsb5mJe+qpL
EES1hGMeOpdvUPLLJe9h/dVtiXUDlnjlsaZclbZPmxHgB06ivAFM+65m6P+y0xOV
SiFA1FBnXknqem0JRxLh1jbCcurnRst4leitANZAm+iSySYgNbSyToM4O2VJippL
vgEO1791QpB6Zw9z3mTp21kUdYnThzroRuPDh10dv2i8KzLcS9uTaJJ0jrInNH5k
NG30J0Ad2F3Cos2pRfk/OTCH08v+qw6Oodrc25YYtRrFnJLj5m87bt73ppAYX4hw
7BH3eHRlaKeeqM6HQYgkFfRIF/W5hW1ByhVYsqajkQmA3R04vDN3l2P5oK+vzYn4
mGdsq4sINoRi6rq6gsYIMyCSlpnov77ZzIqQ1Fobg0P5/ToRg1A4KcKCXVnJpz3Q
r/gmCRPGZ4uA94weTgaCTKPayt01qGHbzEHNUuc6PlJ649wuxqSfj0vGZSqRmqC+
TQEVvUPjsdZGha+2QGHGhBR0+BicMjFwIgmaTTbVohbk4n4USf1J5/MU6zQhFxJy
AtY44/vlpLOCDCf58+/odpaqrw8sT4F/0CDdyqayYvsv1R0Le5dwGV835gNb6s+Z
xH1vHqcy3CnNCfwpww+VBl7gDGod8qUmWkPTKu9bPSrq0r6TEyPJG7CdQHypv4eE
lc7GyPnVaz3CiUqEbPOrVW12k51i8vaANU73GbpNxDSaWbTsXl4c/q9VDkVqlzJ7
A+XNr8zy3EmtY5BiMALoOD4gqZsMUTaArZyWkGwcSVUInKZBvGlceeIkq+zhOX3w
Q8EtspD32GEJPRj3Of8H+OOPvVkh6zYAzilrBWLzrjYaWoImKZFG2iTISSk1EWwE
/vVSO9JAbkFKF3/bffB007BRFvt0o7dbifUkxnKXY6/cEmbnONkda7GVP2lZds/8
QkKP3NDpVOcvN+rSHNWUZf5wNk5g/v8a14yi8N9a6MO0UARzLWS8/IazEzigN9jq
0DZmjWVNz8Wr8c8w1BPoBKutKdZHtdETldWPmm5eEdFof+kPgy8Ug9hVsSFiRjrs
zO9nSC/0l6OTk7O1bTXAtLItmCMkSnU+a/77q020WtpE0cH3okTnr0+Y6ZTyj83U
bhjie7XkP17xnm7TdCXKeamQchbNZQeSUAaqZMSJ1btk5xQPzOwGNfJlkNDFsEcj
CSFSDOWMyoxXaLaCQd/SLgif9DReK5Yvol9/EDnLtYiFPfi/dkjnOSeHQFl0b08L
Il6NM1FcrTSIC6cLVff77PeVJ57djTuv3myigtHTDZ0Ni2X8NLMCHm/ePjg/5/gQ
UZcf9wDvB9B4PtPes3IL5us70Kpfc3GDTHdmUJvlFqyNtdGnjwebyChQtjTD3mks
jVKlDNs1iTidxc8bzxe4/UzSc1rjD1ZTcIkxTx8ABJYC0zuOHdDvgYcc/YOyb/Wf
06Kzsr0YYqyMkbBsBuikAkfMGXMxvYRdrHivpW8gTvJBUi/0CI/eD44E3qgn0h6d
PJXSrLL8A70j2W9hEntn8kIETzs5qIzALOoRIamdwey6Uex31q4UJ2K/AMYj+M79
t5KcHqs2xvgvxTVC28p4kiXQyTaqypbFEkzp8rfX1fGaHvZ4aivb5zAvMkPSjfXk
W2l1ceRYJQyIUPzoNx19M9NiGZ9vfNY02hgBjGuWPH0HC2CCyB4VEBd37j/b9J2M
DCxj1jubGAbTfhJVQcNHY0zq1YGc6Uq9vr5x5TqpTDb5kpBW00p6ONgDCYSOA9HA
2jYusVQ0v83cM4UiJ4jE7yaXECXz4TzDFFx7jSSkLF1XX9y43U5mmlqiXcO/G7Ts
x6Ncn53jVH961jj782kZNDSysutz1qITBlLK0Dt8W/+8FTaAHjssCjejzsRhNBCH
isQI7QUjDFHCC/NFMe+Si9fXkeLxVefTeUV99HsGLWRJh1U3/Er/VlGCWmarnw97
gUqET5Y+IhEffCG06J0E18YuM0YuXNfNLP2R9TixJOcMmaFNcz3Bz2X3KBYMkP8Q
1VmnGowBI4oOpnehqqRc2gkcoU0CdBcitn2pfB8XL0098UGAMuIcsbyHY3K+b5gM
N8YaDSw2OYLusBtGd2HC+390gY5PiFJScpLu3yEdUcLnwPMePeXn82WS6vPct0yK
RQ2QdEgBfaNPvln2HZinwgFSUU+ebE/NR4em24E2PmRJNqUvKMAPqPALWUfuRi+k
mqWyTSIOvDkSP15jy3HFmcqN3CA3z/gguK8rqu/gP1mgXhA+Q/p0AUEDilaUoXn8
ze5v8XLF2vMj1ET8hF2URrDipiPpye0c7CiA7swOKdM5tOZTtZ/PfANCxru0AY0H
+VdO3G2ApB2VzR44u/r2apP6wQCaNX0MoKAUTogN0q+CI3bbTi3IF8O30bsFQUW8
M86rVHEsshbQZ9Aa28ei/isrlQqwQ6NP/Ly6ZWECwQsrh//zSE2VOEm6W2LfSBxK
IePzOYCtrSexHoFIflsDViSOwwjsQBU5hlBrP513w0XTMRSqXAsbC76cEmj9JnoS
YbI3yiexCB0zuegIA5mUnGfUQfZb0A68ELKJe21wn0YhrhEoE38N3c3s4mp57AjR
6e7HE3LVsZ0W8f+S7iubMSq8LaoinZnDSLbPqTDvPirK3mQ1qc7K/hXcG8AS557R
pqHQJnh2vwKwv6VgPDSaPCsULvY+WjXsGDow6Cgzk/LE26ZUnburWEiY3r2N841H
CoOQOS9Kpy0m0ExmZq6kkZcYtiRIwhGNLl+xU34dRe9KJE1c1YH395Zfhe4DIfca
0yxEv/k2mzyabL8tKJmgydURCL03dAhrRLv2k7wpmGlpJxDzWzLglkxsocvL91i/
shjqANk1BqKMOq5RrvJDaazdm9tQtCm5vKidTgkA7Bbu8Zp8P03KGA+7r75oIs6b
huESoSZek6E/l3fz3woG5yeiVU8+RzoqQCX/uziclrL2JcgQ/ddTqlHEXYOePoUy
yG2EtU1uV93aePIxi6qM46KxNtfXw4/HgEzCfxbB78RCSBi0eVpstBKTH7MhS8/5
k9FklY4DvKVer6VdDDDbTBkDHNJJP9jSMwdFaACQglnHxNTWW95+urO72xHAWT5P
aYoJ0tKgbkv+IfBthfE9ja94Vgp+Acis9B7XujJMUJQaPX6jg21oHT14rwutnsjY
t+U2Wl1lWbpUHwA4WEktdcImQJ/LbxnMxEl8b3ZC6BOA3YS5oyQvVwZOo76RV6Qh
gNF8T3OaT8L0DsCxv+dNvjBCTcKvtEifrtvlBbit4iIGeY56t5LzVvTGL5mbBQQV
2kaciRqHA15/uo/sEaMWXCW/ToW7JUms+wUvwdqzbNbHf0pbBqlTITve9T09l6LP
KoYyBtUr5Mg6aFUc5r/czVSF0uHpHD/PZ9Jvt/6O0hvBi20uz2gCPTVC2OWmje+p
PxtR7fBiRZ3c7rA/VE4R9RF4XAhq1c2h2QosoX0qb9meM+UCMMwedQV2g9FHyKVk
gPewj6O4PVzonJB3cfl1O6hPs/IRFepO6SB0AjOAp+pVSn/A/M5qZ+xR4OQjknmu
yFtfgEWbFypxjgmoFRG1HGKx68UVQ+9T6CQikCrgzlo5PFGG07KbpZseOiHnbIO1
m1ixg4j8QJroOS1jCFZMqtJQyvbqV3BW1u/d/5mf2Qbq6Ra4yXbP8VnjRFOeg7gT
f+JG+woFLQ69/LziZ3Mf95hOJTZ8fG3WKk4n+VM04ygWqEHmicz12pAO5+QACK0E
4mv8eYg8SRqjwOzVsyCuW+IVRnr4THTUHCW+Lji/1JX13OadjZVEm5babjWiVNUD
2LCmjLGaTsePoWJTIc4WL9ZzXqQIf/iQp93ylYqlxoTzuplwpdF0qRPlXR/zDv9b
rgXXvdrNx7pnMR/3Nr8tXYaeeDpBosCe6VAw6np5h3OKVU+bnhb76s8wyqtzx1ws
QSx5ZrleN52nrOCNwjc4SuJ4INZ326YfLQ84C7FuChEZhG1/eB6zyWVR1e1izZZW
fCDQ2+YHjF19qIeMppo7J7JQwsqdIA+FcyahxV/4f0J7hvdlwywDjiklbr8/gU3W
kUXDHISgByCzEBUdfohqcQiUlqiW61uOBRWmahzZVG04Cfa+t29GBmRK/CNtXsdF
YUh4e+4oCIE58l7lrKKL5kwZPQDFFm2BhUvivSjynhh0S18xioX893qx0MlgtfQf
+/Z6tgp8ukNOLHi0euq2jUdhNi3WuAeFXQfbfxVuR7swbwBjq4hxVRbY1/15N63E
X2eAkCGZE0lVV4UAEjJk/LoybzCNkB/FJd5t1HVr/JrXgqUJB7whQbCvuF/ZrUdC
rODeEXeg3HrWZqTLDYp2kPM4KA9wAa5hHxNa1c1nHxtJK1WeCUVijAEKuXcMnuOZ
aU0NmjD2sW3Dz1k13HbvsWeXUFy+OF9OHxYK5voIGRdIjfQHvME5T296P8UHjz/n
iJHPZngha6+mm/o2I4f3WeKK08sQAKeco91Yp2k6vWF7gFKG/LTUoie+PU1cKkfS
Tx1Pb2f/YlskR8Mc7ocp2ygOB+aVkvpb4OXj9h5k066F7/TUCdNU2FTPdLLmepK6
oPEUwbiDlX8XBLFAKGq44w4wm54mCUx7UaVvCHBATtjJrKYS4QGdXtKGW5r1I19i
DKbjXpFehwi0m2G2JQ9MiF0MIoq38ZDFu1p8v/Js9dB8spMMGJGmq/DNlrV725Hp
XG1eT7LlFmesR/5NWLu/jlOcLhOjC+cvRKXSQvLiBQYYQiF93CRZ2DnmzT0AIydK
a4RhFm2q1Vvkz2c+20ExOcqhxhqd8Xx7hU9lhKWnKaNQ79JRguFXVt2oQ6ynhtNH
DDhTA7e/8xKt/0RnpwaYCq0Ttp8mJLndYDoztdtndh5NboKUB6yfjSiOT9PDcfzY
Tw6s2+YQMWmE45NJ3oU4B97nLS3dThJUs3a688jagCm01fJj7sis3X/Mei2zODi1
2D8nVFzy0xdhwV3TjoFHei5Bt4vhvLV+d7fr4OM8QNGV1SHCEnAY74XzjwaCsc6l
wa97BCH3JVoRgWkTwkpt2/rPXfcqZkPFW2S/0MSGY5xgJdJTNDdUhqQjQxJnALoM
nSCgQ4glKvauRY9tpDB9m1Xce3PgkjQdS8gNsXN6z0g8j7eKjnZFoP63iAVdHFC/
oGIAfV7izmNftt9QyY0JX6ojKNBarSfds9k9rL8srFmbtumM26neDwEtACPmlA23
GRHQmnGy+R9y/qhBv70+/KU/+7jDv6Wu7YO+203KospE809ZfXo91ABY14rWogRe
02i3KQxgmQB3z8rwtLXFitEZceiRiwHiKFM5lLpjw1cOITAFd0Y6gbIbFm+bGrOC
EXgTh+3X2lBPzavYqFGwc2mpBu02pVe595j59bWY47vLVHqGIj9kQ2MgRer1wFw6
OMwf2toAxEN9X1Cx645jiOg8yLflqv1pGMWbzRDH9W6PDR+qLb8eiAoHCH9sjhdQ
m19AJX+ncYBKPVwpw9/qNWH49JLCwtr3KqMCs0gS+XvP9XbM8efdfFnSEovV+0U6
RyZttbU+AtyIJvMrb5euQs+AG0fi1qVzD+pN7nTg77g+sZnK+WgoZ1FLsjcvcyTA
T4Bsne7jRhVxa01CEAt8a810XJkWjP37M9A95YSk9HMkMlmIm57xK1cWRcy5Ar74
cPpDQqTdY9Ljw349++Nt6cuEORTkF7Nnx+q/L5OCaW/ZRg+2imeFS9TIA5NlWMuX
Bdw84td7ix+fbCAyhvpExvH6czmhS3n9vuyrQDgfd2Ot9wAlOZaINLwbL7sZZyOs
5TTDjlVSkDEB2ks2X0O1mzhla9C+MKuZsAgD+eKXR39/+jX+nM6Axx3RkQhxkVeb
X7USCc6eA85NaVuKJsfIeRCJK+p0FfJSWVJ47co4cf624laDSZ5h0OpKeBD+keik
/fsb4roU+LjomdENNUGz5KDyLf4yp/VFbuKio+MSVm55aa03YW8J9o/tRqbUTY57
f92JVoJ63onbM6raR/Qghbyw2U1hcEgdIVmaTj7T+1nIBVlmPjHVWfROJc2fA9yq
IEZlCfV04koCo7WlLqmMPR3OF2yP1G6065gsYrxRABIEXWuHC95HtXQTj0DLdBAT
AnhcNRioTU2ZwSVYpZZ2Fb56S9761H8/H+SEWORSctpKwV+CJ1CSoAvVYXXp45QQ
tQNUdcEO/N/hb5rhT9FAUa7pX+io45mQBr2KJ0dxd2OuLovz+bWKBhFJ/8Pyr27C
tZKM9UVCtTkeyt7OJQZ4lmd7+D9uhud1OosahVdUjlSaGihqhXWsCfVZbEx7XNfd
T/QOGFq0BknMM63UHyTx89Neljj4Lnugvv1J/Q/F0lbDmONfQjhkH/SykN51eb5i
vFro4Y5ikbRJ7aAK6P4dKnSCAkE0KbjpG4XGCb9H2vfJz/8knb7twIQTaIwHyx4A
djQ//zbv5ZUqS90FPXpQrJrKxzJEldE6mXN1JKc/PZ2nre15ZjVRhhfWr2nnLPyZ
pc5pYEthvjiKiu+u8hruiFGGc0FX0y0ZqZ/6t0uGf5Gt4J2HzirfmZITPYYR8oZN
2hlBhEpv9/iQWeO4RxNZkaKWJoz+itRSuwDrzQYVMjsF4/P5oMshPJbbSW5o4XCa
Ot6pKFqUpvCmxhvuH+3H/B3FdPaxZlgffCJLdCA8h3vTzr02ktYszYwJanNj7yYK
FPXmjratjFGJ4nGZDk8oo8bbC2mb5fsH8BIreCbjLlTm8ksu2HpE5/l3Eeo9Hxcx
Nie8xbJZ4Aje2XRpDkpxng==
`protect END_PROTECTED
