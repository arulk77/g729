`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DZq8a+oxdSGJOyhRMNdtE6IEiMH/zihtH3uVjv+NH60xKB2IOn7O/IsCgHb88K/g
xnLhSsQ3fViKIm/Y0hqShgbjclGKGhp5QsT+d7DjGGoXlLG36J8Bdm/vhlhThoCs
04bsxINcEXDQkOAsyGt/k9Sn6W4OcYIhdDqRXMq0wYw2GaU0AaMOHLS0As99NUBO
efNr/Aa8LL5sWfheq4W4meiEjcEYNJs5+hp2MFXBa6o7fNv5jF07m6O16DOy3euy
nA5Vd7/sqSm1ulCQdpdnZI5WybZv54GkO0RiFCG9gQShKZrgnRcpc/V6jWLeBn+q
idtnHeyHcyB3BnzHNhn+RkPzD15byQZojI/lo9HjOk7uO+HyZju7cAsL0IXHpXHv
O8+tCkyuoFXFEcpc5J+AwV3A+8Uaf8vPtBx1r6GI8QAjeI5fwnXfwmEPPR5DqLFu
9hKgQFGnacOiz2aEbg5Dw7Gpkzv5Fc/ej2YFSlCg+D+rvp/sCMDWVPYR6vr+yPsm
KBGqWnIF4rdiQISMW/dloA==
`protect END_PROTECTED
