`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDkTYeq0UVt6ljwATFp+CmVrL+dhrUsumAoXY5EMenJj
24HoKZ4O0A9NJqKkxu6bIPNKXmY4UhRMQ8x3Pc/vfohABQ90gGzfHg75PojMm2i1
DaJ2PJyerEFr9ThmGY4DJHZxEZ1Kfkua4bghzAoWF16YVtLF+fLkCJWBEU42peye
yikXKcmYRPXrL3Wprmz5Hbp+5nbANcpYiFwd48jnVStdBvcRxgGHSEPOeac4cxtj
4q1mLlH+eK7Lup4DwTFEfMs+x2oYeMUZvTjLf9naCPC0d/eqoN2S6Yp91Tqfjb3H
BUSfOV2IFhRu/dsFODCCJouxZ1sNu1nWo9pOI3lclmfRW11teA/jpXQJJdmnlaVK
xD9w1JNfksr5EpIkB/zXXr4T0vt51w6vTw3yNseK35dtYwcPvxMRlTJYtP86vyoY
blSrewNPWOFe8eT5p/wGQ3Q7LE827UK1NYTJ3OD6UQEC4QosZk8BrmZ3D/ts4Sgs
ePiP5CKpiL/xXUGBkzMisA==
`protect END_PROTECTED
