`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveArBuraDe4fgYy3NxxUSKGgx1Ay/4JCM+4y4eSbM0t0e
7z435J/6IOD0qVtIJgio7nLCGXilWoYYasuPZ1UDVXP8h51giTR+azbFY3KVt1kN
hoHXqMlpTa1c7u/HoSDJSXIpxWrz58LJ5l+6wrpRURzZa6F79rjCiiGf8g2vWCPv
8+DNVSWVlbrBUNesXKbysLgJy748oDRsfLnEuHLJjcteKh8Ivia6lPzWVeltGuGn
nuGB4N8iEm1yn47GgeThOTqJxv+mDkzYKMEuLLzhyZRJxFxijP1byZGY29hwoBh6
o4fau3rIMylLs2ztxcbxgw==
`protect END_PROTECTED
