`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wlxueyD3ooMyHNqibPSHeQ076A4s2CZe16DbyRsoHbe
gd6KD7dEdccmwNqHHWValTBDZmJCu0A8o/+8Rb8rbLf5AuD+qNqJmtAo8SfqqSIF
esLO9AHeWVWnbT9/AHIG+vaF19YNfr7rhxvA0Oy9qNtohWYG8LGlm5uqBWs3uvtl
t1Zgf1huF4mUTOWeFAxl8Cfg9cDCYFhsAm1ASzufAcx4J3abE1/q9tuUkqCZW3mG
ElMVJ1oK8k0ri+1pfDd01jwXMJP8MPxgZgSoggnEcQKjM0/+JtaXoRnI9AafkdRj
ZWK87deK6UFjgUmLmkX0aVVgxXprWeT0xjzieT+w1sO4lzZeF6BFvXT9yBv6bG15
D00/0u42ueHo3MEGzSyxZQ==
`protect END_PROTECTED
