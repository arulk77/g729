`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDATckaAOj7PAM7of7qhNprH6UYlKTW8xB8ZV6tXnI6pUA
EW6N31ZTiLvTq8sMMGp89YZEKElAyN9x2pkIwgfWr7jHxs/jlCvi+hx+l2N/Y0Ut
Z/xJPcadhm7/Zt9U/oUhxIkF1NbPK21oE3ap5Q27aqFGz2nFGAvTltU7WtCLLHMI
NppLIW9CYtDWyYnqswylNUDV8/dgPsFlhjDO6Sj5JZC60jA//IAunJLirt8gKYDj
c1PevIVOHTjGajTY+8818e3n9UWdTAwOXiqcHiY1wlYZjzheUrmxTSdIopWzvEIl
YEjyGjR2hC6w/QJ8zN6JS0CA/Xk12Q9mqTHFzxUIJKLYWEP60uSA/frEEgqTFBjq
zTaRBEdXcxcQD1SORUyMcPYP7wD51qwH1+CnWvz6BaiiVPghLIEl+x/u2BAH2kGQ
vgoCj9FtenmuC0BMbMZ8R9YotJCJoE9cnJCIGbyNxnW/3AEowabpl/S3UIaprECG
ZOW8F1idsPJlD8nvqVnYq5W/hXIivlYKLDMjjyKgTvdx4tITO5Mrcg4zJfCD9P6p
aPmpQa5Z1UvDHIdVcX/9VAm9kbkdUHE0tWHyO0BckYlRZhOsHleYHmDeuOWUSjRF
CdtvJ3xBAfdtTIcB0EkaRU+aCHxEFnFSrH/0q9h77j2Bx4H/oXyLSQ9oaj+3h5Yx
NR9wtDouaV9B0ixT5H/iwAakixfSzyYjire0c8LcoyF8k4Z5rhWRiM6fh9QZz4ms
58/qUfrA95nIxIyy842n6tlZ7uws3nJhjP2yhfR9DZ/iyBTZJG2xyNTjqpMgJ6i4
xi3CrhYvQy3C5CAuCoyHhDg8kpGtp0FC7AXqK0JuihYTwEuKDrgWSM+XGKkbG40c
JM0JBhgHSmugecNhiTQ4hsZBsR5daxcvC4Vra7uoKxVgiOyO/4dF8nd9Zg9IDEyh
yUna3Utw3UHaPIwu89G4NiH82f/SnsPe4SoV/tQw3G/spMERjcvqRuRVqviM5AHs
GRW1wSubhqyI+mgimkWpVakbumCcSO2huNRpUiWzkJNEj8fHM8Kp58P0btjT+n7h
d7txPfo72QCXezDVxvkflXnSC4/5Jcr76XeOcwiLNNvcqr/VSXG/FjCwsC6wiZwZ
2d6H1RSW+wmGEaeQSv408pCbQCXKQ8C5xPY+2+SUhJ+8Se5fZbtHZSij0G9owCYq
WP5b2KsF5FeIEhVdEoPVm+LBG+KFq08gad+SQptbiz3u/7EfqzKjIQ6xnJIz2nPs
cVxFvHBV3Z+hIpcvAgjIJ83y9wlk6PbNJ3e35XLcy0dFLAIvsqIRa5h2w5gJvFJ7
MKCQ2Mo80QMbChmgJz1gNeTcdouJohvgW/HFTBZ8pdxmS4zFDqpUqjmNDNUq6tsS
pReYK8j+QpsPtCWtiLTbG6vwq8oh+AqtubQWkNJiB9uH1etEvrNy4PIFSzOGj1dV
jv9nnoXqscS1P/LMpqESQQI79F37/AGn633riZxem4/M4pAd1kkVxPEoDf0wQtsG
grKrwtjl7Ech+x/VPygE8ojhIsdErkUwfSZJyPGbxuLsi8gLqyxjivQe3Txcs37W
UJfftR4t5nOu182Z36qRF6wH4FXlsx2H5TCbwrvr1TMp6LNld6e7eiQ1L8aU46Sl
NJVmoolWPRpIBP1PJ9Rcn1xCNyu/VpbbCl22+hy5XzHPZ1LW4v36Tys8B3YHg0sx
bDrcUdHByPICYrXXp/a0o229ARpBkNX02xUViuTwheXPTHSLMZXgV/9PKWdDoGNZ
txuHj8zAif+lxaMNW+8EwpIeHcC+EfUTTPtd5oIQtDNHorfHj1/gprz27W4rFtxP
nuYm+nJDnCpMc8ZZPSNNz1VdZEbjGq2U1eeTguab67cg+bD746032HIkgJdalw+a
9UhvVY5aMUl5TuDrbuxFsa8EyJzvGdltyzpkZui17UTqEdB+ioS6WuTKOOVWxZaV
9SXckw69Z8x67MPdBzTyujzwsPWiX0K8iuaQ6WbOH3fpp3yr58pJMWncxEbMFmhf
fYS/ajWJ7BFOZCOMI1Xl7pS5L3KxgGpkJFhIdbWlslegV5wW861NyKi1qeQpcltC
uJj0Q2ZuGlpQrePMjd8PWwSeZt9pd6PWgsLbwrsbqV+Hdyq+Lv34WkR3UwcLXdj/
i71dXfFAyN9Gf+DIKsSiUYMHIvKFcUg3Aayw60FrePndeGnbV+fODWZCpzfpspHE
/J5FXMUvu8j9A0/K1u8CjGp7buN9sXtGOhrxEYesbLuyhoWgbiLjynO3DSRh9wZj
j/ItbNfCVAXjVsnMR9xSYoSzEwQ3jPjKxmCmEN7gLfplZl5Ix3/ZRGGAZ6I6n/KX
VI3sz8hRZWfoGVcD9OLA7XGKZMBKFgEXWKvx5NmQOqrUo4+y8COhV+xAQOuHp9AK
4yhLNsnEClE5V9ZnbTKq0ibHGdlXSr1RG+yn4GlZ1Iq6V72D29eofa0jphYi6WTs
vMIpSqhWBk7mKg+9TbSJ7ih/is+316NjiB2V95uepQG4EaygELCAgKz9Pq0Ecrln
25BhD3IVpjXYlDlShZqCSw9nEd2na2wetqwwsyy9M1gt1C6TTHvwgwcLTp973/6b
8F9UwMi8ULmhMhvA1dL25RnlbfoNAqZEDcQLEgNcU+cWt3zxSXwXqkoMHjNHrgWs
IkJlIKM+ui7m23KkSrmOnEZo0VzalRUEkTzKgOMFI9E/RU92L8RoRnDYJgEoQwkA
089QGhdNdt+0TLC5Ar3VCFjMo0wiKBizt6ngUCn6A1uueszvNguYQI8WQWk3pFwh
AIU+wIrBDzxYLftbnBJb/paoMP/uB/AfTuPl4hQfRY5Lul2AlRqDshedHdfHhO05
HHkRFKvOh+mzNL2MnRk3LLv+ygQKQOOmahxYx0RbBcDjMZXkT4WJVMrYb3N5bwFZ
sgB8ndZDqz8lWcf1wZIe7eAtfqDsa+Np2/+wQMMat3CC8F7hNZjY3UbX6urBFFps
T2mSQHqisaLpZBysGyTDNoSIu8BeWlJa0iGYDImkqUl0V+RZvLd82A9gD/gY5ohh
8XJ99NNPBp+BHJGYkUsKx6xLjgjGF9b2cxvNlc1M8xYUV/V9xtzA0oQTtIAB9yJj
B8plYsJRWrTJAMLQKTLtHujDK8xOEtEgnzI4bjF6JMaL1ms4OEI/hdlc+9kN1Nj1
qZo87nnOshlSwPm7iqrMdddeUHINAFmAI0eXYjazjcdiEv21SIcU6hd4/AGTuzJ5
SkxtqziCoQ4WytftFmnQGN+eEpV4MCQzL1kh4rynigCq8xA8WbDkGbYhbvW9fGmA
z90gRi0ad52rj2lVoXeOzRoqWY0eaFFcvFWq1QCLgRKNUngkANhwl1/OdcaYIIIC
/vDjb6NrMarifROKMuOxiv8eBcFHojz680IQ80bp4Empi5/gfzQ3aNoxuPBQ66TV
gAxftwG3V098lB3btFDvavwtdKCnQsW7QhBHbT7CkF9P8zFRNUvRK72Tdyl3Q8lF
NINEc5acY60RNku5LLjgEegD3k58r8g6Ww2WixRZjBpOeACFeZ58G6GZQksCbyUM
4WzqIT1rtS82i31ZjWl5asIUpyjaeWl4eNbP9S7bm2TNpiOpAt4TXn8eWlREt6hQ
OwVm4h3gQVGeuJtbWrhuT7fkhGQEQ2PHdKmURTg5Vth/cLZcYHiBBqG5Tx6oXXh9
tVFjyWjhkESrDeHl2BAhLO+Q/OEFyrShnYA7g5qcq4wPPfPOvJohawqCXxqIVsV9
xqqoa4gU6+dcUgkIzhyvBdmVRBw4hZoP7bkQ8MJSk1gL0E0LMWUNY/otFah4rCES
13jMDAJFCBUC/e1TFq0u6fzXDIPbMJ8anqaHzskX4yq/6yKWsJzI35pSfmuxVUNL
OVfqOjNCNmVxq1jMlAK9lCTfvgyy0mT4GFvIKNRLG/Qc30SrY3Y+8wMJYMmKKw4T
J5qBFh2/3PLgKgRrRqZVFqnrIjGICLj1z+48Q3veer1fdyA7UE6JLP7+TyJrHWzm
wRWMpGizeS1/B7/qItq50T3knWCTfgtq0x0ttka32N2P7QQ093DaZigAA8MkS9Ab
PMeLg1WXS85MRke138066n7E6n+erzMIeZI4qCFEhjC2drA56jES8yywxTScQ1ry
FxtukX7f/86MwNJ22nK+F9a4qK6p2oD3DsdnFU1uaEOD0B019VNwKp6GYpLOExmg
psORB7v3a+aXlsd5oc/ZHbNPXy+lIFop/gu5VvFi5J5YthGu/QUksMsgeTcC18mr
gSYOomI0E+iUrBDTBSJL36GtAKvcwocf6aKDjwyFQXz0r0L8jZHGTKDcSA2PMCGR
PpGpY9k1zG/KT4UwNtCM9S5d1wUMh8vaiQq/thTVJKk9tnnnFZRiHIVeD4Q11ywe
UWMMlDHOvL8OLuIlLG86ywN1zE46ALrNH0yU7FOxK9r5avawP037hL/urcza+Ct6
0Bgt/+2btaWndPStZ03wWTUU3u9yP0P6hbx9bMPYXLOExkMbjbLovC1cJEFSBSo6
439simPHWoHcTIUJnN5x7rMckhhB5E+SPYS+H3F1ZYucn0WJFnZURztW3xaz8OKe
RvBj3MGUaQTVfgzD5XcHPNnvH3NI2IdZFD4Iq11mCjVbSUuhK88O/02ewXYXdhgZ
Mz8oKRPMzahwFrvIwSQZsWDxNzfhgIVPPLPDUCOfSgncOZHLfXQggWMsFT0/NFl3
/37Fkk8A/e3k8NIOlqmftBEKeap2LX5QB1iHzswLmhByIaGQG+XtDKtCJYh/aESv
eCuKThXvxMtpbU4KcTIjYaUEoPyX0kehCJ7as+2+wwX2pIOyamfhi+sneysbI3up
CpOWRgci+/T4XQst9uK7EFpSgqCfeILhAt53x9X2YnO84zLPDedOmBWcY1LpTiVW
QVp3ogOBoGOeeSkHwEdvX3Y2K5I9kpWt/jwn/oucpBaIzoCDzmKz/tfojKAdZ39P
SS/s6vXn/FKpiiu/oLA9/mhPQOsQa1AopO0+8iOcS8UytcI8/Y4F6Fje1iilnnoB
key7YXd+tQ1JIskv+ITzE4schwzvaWknALpNpJ5Ph5TUoc9bXWOax96kOoKSBI6g
qeivJOJ/x7SVDqtpce6OD+d0hB8PxYRyYKS56WaItQzgDbWwdRITKGo3k7J5McXh
jx8hgeu5KDuVC3AMj/eHxLIWh9+wBPvoo7WRK/RUvxLi8e27zsdT2/DbsNipzzLR
+sOOS9zsqZiq+M6mqCBX4qEJoVh5yomsNVKey44f4r4CbpxxIZSsnXCc3+rjWr8A
iqCIf28vUU6P8Bx100zLBXsc/mbTEWac9Voh7PN3T987aHo3BWUcNSuNnCg4RKIv
y1VaKZvPuTTIC5+1kcya3aTGYJpxcqesB5sufCu2tQOrt60MKmKbd+aBdyRskbGA
HLMvgJwqlkvGgXvK4nkhnWn2Iixo1KfYQi8QWJDJJRJzVzVKZIw4KbcH8Xmd7RSP
VZh8S7K4YZC82GRIhB8YyTRE0HNgbeMXuGJQw9+7/9aPK6qxyTzv0xQYhnJfphzZ
uljoOrUfxuzoPS7u87HZiBnbwtkDtSIUrwU92nRdU3b18Ts+7+8UATlLmlp2gVX1
b3p2dmmK67vWdd/JlDkcPnN5fKe1TOUcGrN31ysewuLEdhGdYLcOjllmObmU4S9F
gZ2EgSXTua2I2z3U2Moskn7EghIkcOTQkPYcwRe2KzEzrGhr8EsfMtp1hmjIHxMZ
RVP1XYvQX7+w20CoggsC4PuBMHi5MWEKfNQTJGC3GVbLBlMIpPw/O2Af3nijfMQZ
Wo6xK7LMfgjgaM2fyr44MEmk4H5cDvhH/X4V58nD1RU4dbnxlvbNoxCzDHKU6KkM
gfJO3EIA6FFlId1JChxZlkSUy/h50jWR7SdmgoFsSvfKciet/2/d4fWfGwHkHspl
fZnY2koAJD/6y8ipU8MH38xzfdJdkcntegxMatIyVigM9KzYEhxa21tmiQbBecdU
eszvD8vbQAZOl87VfUkghkvUntahD4597mdKs45uoDbhbjrdB9b6cDYlYO3XysOl
aFcQ1sdcImRYh2A5JyNO+azuuxU817S/df59LWTbyPwgD0nf4zRetK4+EHAFveoA
69alnASnuLzHP2NTufrkm0/2vMe3dIauEUOfhykoidW31c2EYzn6vBCvXP2Eegth
VLNp2hubiKcnTroNom/rjCp65sp01pWWyL1XEDlSlxNDemw2TLKFsCILlPfhPpwY
K7Q7eF/VhSIDva6VByUT0jLQ6OQ3ZiqTrTMbUZtQKIvcpSpuh+8H9bxxYewadEZ9
2jKsQiCDdRtVR3qQarNNiw+FZF1KsKkpL7+/BcmTIdxkQR7w57IiTGQZMsIR3FaN
Ctgi0nXZRfPG2OwgoFumzYO/zg21lBnWaUtTdkLFH4Dv4/xuoJVSCo2OpZ2bSNix
pvECWKHBfxdjryX/D8P/A1ScATbvuurybEBI5cCplxKbBU48D0GyXhTiCOm3UkmK
hhXaDD1ZbL2Ee82SMGReywIgFd9CQKyzSFTcTknAL3bCp2ySZ6aywYEmYH+kfpnw
AYXSPkfYxCE2h1oII9KkIerk5NwqFbumFvNBAaImwjTHaP23LAp8/7oyCXd6eaJF
cgXRoU/SgQsVOrQntoy89j5zu5vBSiXcVEbrur47zv0pSYuyWpW+zcPHzQZKsSQU
qkSw5ySX+/ulNWMa7mut+P/NWXInz6xF8tzzgoQX9dzaLshHJ3vm0/lspyiFJEOA
k6SLBdbRVxNh6xF0CfJFICD8BxNOw8rrPhUKpdZ0osFvmvZujp41BGDGH0x6nfPD
DyqZ8DZx7Y0M1763SRfXM88oRkL86/8iooM8QKI09Us7N8xiI/23RmBNlzUsueuh
Rxc8VaNQj1+52+Xa66uhGCXSTg0DqoOrmpTGzreOM3hSox+ixcnrcvcVmTKPYBKu
TtM4j/j+WU6tLNy7dISQd234Aj8fHixdm6mhyz92ki2do/wSE+xP5GURqZHa8+su
MKx8ru6uBG5/1c99IV4q68+6wR5e5Um6453d0/iq5P7EUsVnP/JobYcmnTO2Mo3C
pA5HChLOcxP1xvCoQvcrbucWdA8jlzlnGOgCk+VQunE24IhkZurFD3D36zaFyo0H
vRf2lnOnHK1cvFbI503rz6C1oUgzrZ4bWwimNGelqHxCnLV/yl9MkoxrmaSskgGg
M8BHO72UvQA3GGk7iPC5yyST/Gd6DnE07RlGeVW0VDjWX8Srucc3cCY2pmlS8MHu
HH9GdtN/2L72VtUbX4Dt0PwFvjA4s5MPueuKj5Q3EKWmTavk0J03w6QV+PcwpnWE
PI564WmUWYbMLNek79pJiY+lgLtl9Ew6m0+fn7c27ffupovuQA5B+BFJ/visLVfE
t/c3hHqpY1TeS4gvIffPmWHzHOZTcj7Ca19y+wnVgV0iv+sAeqYxeK7aGlCPNxQ2
WeYephwSURb0K5KR2MfkDRt7loCXbRLoUceYIqHsqR26iQO0FAF263WKJvdHNjrq
tqhFH/NE92ubyyZNjHMxss7YamIMwmPe8chylJxh6TNCTyixwtz7DdIY5iu28D9+
X+TWSKslnws87iGg4scJBXlrlgAzrnar0qpjysSQhKgbg/gumDoqhR90AIOlxO3N
HfNqjq+O0pBIBzzbrCnmXPrJQFOUyekzT25Qpea1+JEGc0N0J8e5lQwLsqyTerm/
TXg8s8boIBnwTO42lcy2V8m/f7StBYN6hj7GBgewlDo3sPYZfX3j9N8DkZFpYg5Q
PatN7XurysICfV9anBdSnZxrIyGMk4tNhRx31G3WnfTY58IHUAoybroLC60uJT56
/xASgZEk9ppGrpnqaQD0KtI1Tt2loydOTvUvvIAotFk1VCIaiA2YhP9R6yfJ+zLG
bvRqRMXdSkPl39jQummb1YgXMwFTfI6CUZ7Z/wN1C6/ZYkGqyx+349NA8/P780JE
E5w6uvWbkVCWiJJHkdRCW52ac3iO8/ohhBJUk76NmN0KnaN7Hdz5Y/y8/PCidFP7
x1Qo9xU9MtfpAPLfmslnSxjJnBGvyGH80dv0zBAaBZT1by9kNkPaVXaUTUKRPOAF
Zrdsh5pnm2F+n+DoLTP6MQdPd6gpt4xcvBEN+b37Qkm9yf0JcE0Zq614l2SxP6Um
rLQLehyRKHrSgPpSfSCobKGEfjU8U5I0GQf54ZoFuDH2DeCMjc/V3uNghGHMNK+G
cuhJ+lP/uMlpXVdaVlNbStNIAQZtX19cJdSDDRkW/Wayapo7UShz+5r7kfh7plO0
bMui561tObTejqUEyE4+65HB1Jw9iP+VWdxri98GQvGu7+I+RcGyxfKIUuVDfdu5
HVrD1mKX4PGiLBIy5Ao9pmLGPuJnSVA9qc6t0eiu9i3RUjwB6u8XPQKv1gxR2Ksj
e/nIynuYK3sGMKsQf4C6qJfoSpNvbbji2Ak+1W8xTOn5Ds8DYppZbTK7S8efZ/GS
1EDfSbHd0quyofFg88mIFut6/xCP6RfJ97igNaP/mw9khucZgeKaQlXWaYfQ5tR8
Ev9R7OjXGDZAUaGnTI2UTofaVT/jbxuD7cxC6aZ0G9uBAoa6dTD7v6ZYnNW+DWC4
j773GRJTpYSS+7NP1zqIAMvyKPwlTMtHjDX/6DhvRcqLa78VeH93uoCI4cdEx770
wLRiFkcs809LegOIP8kfrWndhElgEPzvny5rFdlicLVPVJTiobL5RgpV85t2t0MM
9da6PmQiCVPPhqBFyDpjN+zIuyXhshPK3hgE/w53VEGqrs0ZV9VErxkloThOwFvi
TqJJFm9n5iG4u4mNA6RGvPpq6QikakBvLN1YuBqyQctpmAuUQlznQnDFjHRgTRJ+
yYXtAenNXnoTL+bAMNVIwuvz5b8wRe1oxbhY3FJpPAqzFXanLdlE50d0MVPzwdEL
U/u+Ai4XsjP6DyDZvYa0NKpAKtwduV431c9ooVae/mce8nnFwHtO8ZkBOAepA8Pz
m9lUBIktqTWlkyEKIySyAdEoOeXE6J5RSkA7X7bxZtCrQ+/zK5YpKzxLA6k5m8oH
3yltCh3lOKhS4BwLCO9lpMrIENbXBodcQfsCYU/Mpyrp2rTuIotwgvDX1/7y2X5F
jDMT4bwtjA1bsOULfvGFBlc0Zzi4B9/uj2nrN0WcUQbDRqZUyiyP2gaKow8CbzJU
dq061aZq5xOP+GTr/nYEXotAGg8JD5C6VIeWi4xx8ObCBidRdvDCkN107OhH7zJy
MvGhZl/sX0khgPLLrcTQoYHoiUPK9cHiZ/b0r5rBr/ssTUaS15yVtd/DZicWy0op
UVuIRN10ToeT+B4oQeEDNumfCPIkZNA4geASpS+7i6XMYNJdnvUnqy5MKxrWTQdS
TNgC4FS/MZqLyx2Md5kVGpbmUl1MmwqLNpLyLK5eBmqZDGjgd8g6viXk2Sf1RrH/
kY7z6AlST1xUIZN3WP5NyOqSPjm1dRcLY1dZK7QzLhJPz7EjHBa/D/mwMfTQfpZq
hboz3vTPWpU/b1nNtRn0ImOLvjENHj221t5vRWv93qJVrXW+88i+U3l8QJ2iHcEi
VGZJ4BXxFz6zJnrkayhHyD16jdQ30V7QujLMnXCp8GHQK8QDHxwuG8T076RWB0XP
6VEir9xRkqo9EYyr95ytmEITfhErGd5TsbyVpBaNhC2ODFWsa1gQkbu1xkUbquie
Hv+LQ6rwopkLWjr9a1g/qYvSFPlV0A8BYK6CR+u2oePEC/jZW9mNjmV4C45HZ6Y+
zTbasT4aBnWY5hnElU+iRWZX/vrrejNI7oPfAxejxHXO+uHT0HzmxQ8gKXaCf04X
i34RWL/oLdET6nprkRFOAxHZ9Y216jMbxynBu0UITV9C3W8i1Dg93aaMvfTy+Jhs
sc/NwBwPI18MhI+dIfWAk525/RIynbzcVziXpXugRJTZT+sSye5POAaNIOZW2YwD
OWojE5nS4M6u7Tvubfl1jtMf7NBgdMx+9AxdsKXKniPD6YfIanxATuaYLCEzj+w/
lcvhX8M9U8vj73MDNJVP6XDdbaFHla0o+UmEFfFCgqUOQqtOR8tms922D30VRuXU
MaZx3j0t6OAZrF4lIk0fQEVgjFFb5bbpWjOhPl6lLVs6vLXOmCQB5Xf1BkRpc/S6
Veurz1oukIOqMtHJgLyo6ydc9fZh4xoyaPalIWxMi8pqjqVKF/ogevyTh2Hs5aTp
Q/wvnl3tPj0PEkCXQMXj37X3kxDC7RZDDCROuXiLyg4TQHNn3c4vcGqqFmuOU/8H
nI9Y1PFWos0Kq8pEaNmLnukQMn3LhwLHwx4PbnzJ6EG/Xmu5K4CWls0Ql3YA1gS2
P1mf/02qzrnFIUDkWx2g2nJxl3mAQ6h6eswG5N2+5DteDKwoRMnJrN8uktcnIgCl
vH6XuZgPL8JSBQ2m3Y6OllP9OE6EFOYe25m+t98PUTsfwDXQReLEqXb35DRG22+3
YhKhKNq44cm7CE3JIbSUJ+ISKXLu43q2L4cSYMuizxst3dH4oSjNE1AIpOyn97dq
BhHbRGS/kLD2qbp80YhQ/s/Hpd6IT2EPScHNnVs+rpsnDMramppQC2ydhCXVsy4k
TuBYffDu4WItk3zMtYGTRNJMMR9JGMTJ28vsE06kw3emQN+O46GV6Yy3NxvNp6TP
aWwGHkoSgrJ0D0Xcgk5F/ooNZ2Qxb8JMzvoS9ekLvLeTmdxTfPmTL7JTt0u5USXP
cDjNq3N3QX/FJARrQeYc/evxbzbjjAsWvTe4fP0WMue0uEvJm6H1D0C6eGXW1bAH
jAgx9xBqyyTtyNwb/y1VIVIgyGAtw3ZCvojboFsG2PY/syCK+x2lJELtRHDxSCmO
76OJt3edC4bNIpafqASHVL26gIt7Fh/3KI2JXYcQifxnC6vAujvKWFMNeangoNvo
opZFKsVmRn0KXYILboxxaT31zCqri90NHjIekpy3P7aeZ8PMppn3vEDbtPi2Biqu
s2FhObl1jqjOokWsMLm1NtxzedMtlvheeFzsIU0qtsXQZgNfC1Y72yu/xrbUzM9a
taJjvNWxQSDm7JHBaIo7D+RPNiQ155FDirmCXIg5B3HV7hagOlMXH+h6d9GB6tNU
rxeDWax1TK3PgGsNZfzh+8fEqdgpNKSp2Ik1JlD9luwCdGVzkIG4Kjt0qUTMcvZZ
3KXa08rf1uMp/zI/ulf65bnKf/QWyyVHIH4Oi4Pz90k9m0yYO2yXAxyENCo/JNP/
vOZAM31WotTJi7H2C63qQ32JUEvteiDTJc0k3epKN4xFSQrDcYC7SfpADfY29PYA
vA0ZgzCjv1DPsxr0xySMCXC2p6Z/zNSDI4vqFNKPYqxC/De3V6N6rbYAyqIWgr4+
foQY0leiGqhu8fgVB2HA5bDbha020CsK4NSsdoZXhF2vBIBXLcWgGBazrCiERhRj
88I0yrAA7VrxEnpnKmS+Rh27o0fvyL+7cLFCyWLdkFNKdwWo4lLCG2CHC3kZTMGI
F6Ra4Nje5ULcb4ld9dTwo/EhSi3wUwd1D570go7Wf7DXtSbDlKgqAy1NkwU1isO+
lEWFnELqSyLMjs41POUAvmhomF/n/mNXXVLWUHQD9Dr+lCIlWgb3HjSDaNFS8vmH
EEq9rgXasPUNeHZ9FOJ7XF3qkkDvHT6eD4JimcCDBWaMpllzRCqQbQT4a1B2NuUI
CpsGNCRjBhwiaTqQVR1ra0UpkI61lkE/1FWTR4LF7kpBHf0+2plyDz5axJOGtUIw
uqRLsE3rnch73xj/M3W2Kfqn6GRK83P1d5xwIOxAbgecB0V2FkbhbFmR12dwQF7v
dBCP2F+CPi1Zy4qnOy27G3jRxxS7XduqVOAhviZrL+cqwrKGe0CeFRmV/WDzQGrg
5TLFRLn6HVF7QwqpG2iIiXVUH8STjDFcUf6wfwKO188LinenSXSXUs1H62pNlC7u
CDg0EXAo4wcZDsLc/8GHJeMC9uBbKHn65m8Xdz5IAJWxfl3B/1DChsZj0wZCdn9L
hfBxXMK++a0ThNZ3ioqDih9Abb2bO5tZUO2KwIOxXnV4xlZXc8Qx0IclMoA09TvX
XlZ6lY6215JIQiRzr3PeH5zVUpV5zXme9fzmSDbWtOKd6NF18Xr2H4UgP/c5Llh2
1xQyScV4NPBpOtSwa+VF8JQsAQ+W8I1/t6NoiBUIXRJTJLF11lflM5zA4uQWfuHK
1hqxqpHanyJD3KwWvnaVeG4xwZDybtH62DIIX/amtuoPwXDS+yudoAcPmKVs3eHL
6H5jU/yJGJXGfZMi6WZ0ENf7ks7bsOyDRIzNw0Z5s/87/HDpuVERcTX9vqwL8rzI
axSKGU9Sg6ZCQ0hT5/2Pam9fmXAnuOIxm5kL3zWa4fK5MSvZ4p7pkgSR9bSKpPdu
FfS192GCq6iQ4PK19ocV+8suHxmR5kN9FLAxITNevPhwTRCw9W+879af06GVpy/q
YvzwCkqDVwb+DyLK5ckxoPzAkSt9/4/kON4px0jjFu3YTiS4eXsCuWaHrT5a0nyt
zlHUnf/JJHhT7XDzpxx3oBH+AdRXbjnXFrUZAAPRVeobZNKyRT75OBc96MOhXCwK
4Khw0k+vm1N96NcJrWC4Q1HP2bmqaugk1dwkGOe2VK28JDZk0XoMiVa1U2XY6pOc
iQjjEW+EQUvh5+ClZw05uXGCJOewszGAuAOUupBotWEPKBT6YShEC1Iuq08pCwVO
a2lyjCI6I5nolIvaO/MKUnspcCPmN49maGw19VjjJZD5dgn8gl8Q8xb7PBCUhT4V
vMhoyeEYGqvpOhVN1OQmvBwbeF8JHmvTtwI0jGXa3CuHZJ1jjCWoHdvvHU785s2/
1mo6JzdMGNcVjLLpVe6QSrCtVwLlYeRlVnFGjRM2uE1NcAuzcdDsnSFK8SSOoTeR
3QfB/XZdDZl67jclD/IddIxX4vW8yOihK8VWviFOMjeruFdYYHojJQ1mlJA+zqJy
DTR3gyfEnOrpnGSDWm/lpBbxx3hFlZ8RnDIKgIIu1jQyHDPRCEalWmOJgtfn3f9e
4s3IJSoTfKq6JbuNyeAPRRxmJAOfQkS9yewzS1UMkvid3zosbt9A9dR9IY2WncT0
bxA5TauPuczTisjJo3qK8v5Bcjg74Hynu9Jaa9/eXTaGCKMRqMAYQTP+bzfv6NF+
4q1zWNDkEoW5/5Yt63mtluxtQ9lQ34cth/k7EOeB2S6qOaExlpMi5sKaNFORqJqo
S7mWEW8VuZTNScCCV3KPhj6OJ97y3DuSr+OZqZ3GVCSn8z9TYbkNfcG8kssKEs7/
n6XuyiDA2HZbJRGbvXRZCLvDgor3unwYWimlylqazZ/Mrro7ElZ7iOBQ2AwK86X8
BV4QKV1SwL2nBK2+vg7YgTGfSBefhgOH29MYDExBcIDpF1V6+64YiOIXLtlnSgbM
KoMLfoRevXKuyjDnJ0zrKI6UJ2X9A0FI02jaaOAky8gvvy+OiEODp7lFSL/hH+HY
BqWcAFRYth+FoN5JV298jPEviIRNA89MyZdOmXTWXKgO4LQGvWLdGF8XN/KnL5lH
BSf950OZZyms6XTdH3J3qcoES0b7rDMQH/l1jQCH6shJcu5K7LvSgJRe66NHje/N
H+lxby78XaX/8gW/6MdWpktUhzpjrwDyE/vWZ3Id/OcmqEkq4PXREyeA89kEf1DF
qBXONHJ3MxFy1GLfqGoUdmFE4lBonozCp7ZMjil9PpzDcnqdMOEPCurIpJC0W1Uu
BU/mDWmS1KyAZU3QqS0IUQGrHdVmcTD6tV0yFy8JUO+cxobIW7aPHH8ntrFRUH21
8Tz2K/93hUoo5/QNq5wAlBEXhFk/p9ZowJsD3N+dD9rgUksi4zRdCl8w5MMZjC9Q
TRyteJ/SOx6Ff+N3Dp2M6Rv0+HJT0ZIoj0iVRaF1Dzc2H2SzjQNnjwGRuTelQbmL
Ivm+2kiiUfENEy4jFUuM/hWzpyRBnJ92IWlsc8IB/lqCFqAGDK2lhI8+2syqkd9q
izdIJEdOiRERhc3+Kgku4jnltDVOdJMHwOG6GNiawNRuRUiWO5ThUuIO5xdwxvQv
4uM3buQ4xwxbY8kXQoLwhQ80xmDfRKthvrvlqx2UmCBeqFVepvRVI+grq4m36lXS
1hnt3/JXUVtv+WZvpgBHdBi5BjElWPqKJfMV8ljZrB5kfp0jXg7znon+eWHgQ1pG
g6i+Hm5y1u4n8fWVnTi+TQYWtl+aaUA0b5fWnDfas7OL/jlG75qBDRqkujBruzLL
y0XXOHl/sWIZIKUfOsw4ezj0GyevPBlZNC8LSmTrWEx5reoktpEomOx+B1KWXa0e
AURhHLrLAGcMajSU8uioZMyBlBaIfK3DxgIwFPN1tRLEgHQLj8IUf6qkA5VW2T9l
nfVb1EzCU9ue2ad7xlATGCsRvnHFXgt+LwMHExDOLf5iZj74jrMO9dTAEPt610EQ
g2jJkvQBxMKiSbHmDysMZf5/JC4konFOVA1DlNrYi2ZutoPYry7NDxqHqxsQr+ow
d2kRveeBDF8ZEZnMW9daDN5loMx7kYmdGPJF6TVTJyF629MCZSytNKA0cWi7nuuL
7piiJcmCO6AcyvLYDLIOeERThKQNu3ioHgzpvD1mG3IAbuQWLWjAqRJfKgf/7Y8i
BaTQXvyB1r4SFrSIlwXqWouPASogIRI+2VcpD7gYlvm8P7u5ryg7KOMkZBwTxK+T
YzA7Peyv54dqeMLuHb4zRTEhCDm6dSkqH7DV4tpAPvuPxlJbYQ8FZm62EB2qrGyh
cbc5YA9ObOpWzvY8emb167NQ6thkBo0c5aaZDKrHQcV2CEtv0QII/3W5/+YTUdhc
Wu3A+fk97rBVghSjaqtcysH6/+2iLnVgpBQzLWmDtHGy6w+icFuwSm75Jo40DAwj
b8veoiiwxlw702BjkFNDmU1yQxAltlqH0YLLmBjLfpoPsMBgHFjm5LLG14BcwprG
EKYd8Q5tvGIoiO0EJmTQYtvsu1AOZ1ISYe5PzfGQlw8A+D+GsqS1znm6BirMbMgG
fsu7v4zhD9h8hRdBvQiyuNzL9EvIQsf6rB0afYWJ715rv1VztFRghPqMD4yhizNg
fgFcPO0MtCv+BAIdTXrIf7HvU1+RRSkp7O76RgIsugs/AFY+nWaJwQVFtQBM5J2e
tMPTUTscNOrwdFnFW4zdSPmeZy5PQSt0l8pA80K/HOCmmPOli4YtJQx8EbA1bbNj
w6Pnlg2nPbubsqIVQzZTzSnccXWd0hhYpLIaguoKVHHuPHuWUiPVHB2oZC9iVTqz
SuaD9SCPRqDLly73ziTovcPmZ90ksmaS+nPMxfOe68r7hWz9lgQVm4DNJ2EiSbmP
HD90NRlpZ2lqOu8KWYwVMNaloeVhxemyJzxs/zeiFng5+24eMEuXFJpY2xNgmR4e
8x3wy6aQno8v8splQncnLZjOPwHitnK9URQwBcP9rkCN2gv74ClyXOvnaRZhSE4T
ymv2qxDhdfdl6Gm5Vb6fqV7xhjoWoZnzBs0HUkU36nURlR2f9/Qbs42Q5ebGNgAz
1lu1NBgztallkfiGg9OvVwiYzY2HNr84JFXmwksuRv0rfY7ZLwLIg06FHfaQ9qpp
38ITYCMy0L0ZksgMLr7Wc2lIXar0D5lh3+sLp5KkqeJ36A9LyF9uNoyw6d0T8osi
yhsO4n9lKyTjRQyeIKA6uwmmKKhpX/hSKVBy+SPQL8p2Ow0zcEhUIMdAtFAh7P7X
ray46NTnWW2qWv/L/KvLtPTcSnBk49lnWtjl+a/IcqPbzGAABvdJXI4OBSdtD09t
wt+5YFSfe48vqbfAGfbFXXNZJGWAvlH3WSGvWhErFa1wHGONo4h5IswDAE8XIY8d
PGHxyDq9KDWy+nD/c2SsUBfWLi88aEJRbRUhwYTOeJKiGCi42zx4X59BiVa3FBsf
9pxr3J7WOJOJIIjBnzZK66sJLILrDHZbLLn+L0SHwaRNuGD1NicouIPcIg4wKxH2
BIg4YsOYn1bCJmxLDNdQ/PTtX1y0JJ/ewufxMhxyvr8fRrKoZ9PBUTr69QFRzik7
xCh1vWBEbmFMUxyX9cgqg4AmrOfSkKwCaSvPaSU/ayKIGmtMR7kt7au1Yvvra4bE
sm4sKbgDqAxBJDY8o/PUux72WR+onvT+7fJtVJKlq4pGVuTAnQ581Jr/avemwDWK
58wv7Ykh3y1Yg5FHw1AjBgGvZtanSEW0U77kb7YAcRsaAm4WjjVqQFYaRJaPw1pZ
m3+z8wJglVUxyRYExA8kQ4yVqg9eURyDb0/Gq7tUTljTGuysVd/dhHjf/vjpASfT
NTDPv+i8YD0khCmVoCYhQ1S4xlUzCPhA5u3WJLP+pPXshVXXLBy5x5QWi9PUZ4Vd
8MQofjGgdieeY+Wml9J8oT/6KEJQKfsaPIjB/RT+C1LeUXFFMTXH6RQTdT3OAdVg
RYgE5tywTRPsZvpqKkcHe//qMjq5FJQuGQpF8VOS95aZ/9l56rA3kPAIbUTLVu3w
V4bkqXr5wGfbe7OVPP4KyuAbujgx9hsjfv1OzvAaMztkHm/b5cegADIBLLXsWN0U
oQ3u9LEJcCEh1urxosbdxpHZdLjoRGk78bEO2jA2dn0lBAGU9nvaVujqFIvIclf9
S2IwmP9cBwiJEY5LycpJ8JqD7pn13L9x82gq2lJiBEgPEqkd3ATjEP9jclwAy9in
Kzd83yOAVKiNwJsjujf6lNJZx9pw6AGExkEcf9yLNmzwwvdzrQQTrPhR2rlgqPbg
PlZJhEL+53vnncTJDfyjxt1XWjBNBPnoLEu9t5ipOePfrDJD+zC9FyoRpYhqO2Zk
96c1FYkYbND4M2fsg2a17ds5HRQXzkjYtBzcHxDIiWLnrfD0PQO6WB+0pkyEfpmi
0mQ7dRliMaX+2R6q6VMlBO2pGrnZcif9x+U2hUifaPGgZ0Bb8/+SsdZIFFp8suAl
eg9N9PiKxQSi76mV01M8lURm3yMSYqmzd/bvOfKZRjm+7o+7VGPZwJFn8bFLl3+i
N6Z/Tdzbga6oadpcpk9Di1Reu423h6R9cgLXoYtkzTUu4EUh/NtQ69rMIY1AfK4h
ASQ/Q/yGgtFd82YScgYXCWx9hmuvQingjthCbLx52/Ee2Ep/o+UDJ1iJZXO2sLOb
IXavdzEvCnByuzlxgfFS+z77dMszrzrPlFDjKvenzkIck98rhHZD+elABFgyHQ06
akzsSWJwzMLa8UaP9IkDkn5dcVpTdB24nOGjCo5JxVR9CjZMlrPyt4/DD0KfIQKF
19YUisyQ5XVvNxTe/oGA1prgQPz9Rnq15aSF+h0oCAipMXJOwnhOjgiUOBb77bhz
an3f7SQo0vX4TonhEVYYJvSoRfSvcf4pe9S/Eg+4cLMN+5Q8O0E+jg8OBFc5nWFk
Ot6huCTSABVZvElG36bOXh66pi/XtlxLdaGWP1bDu3XCF+2gNM16AAfkMgcEwJm9
dhOSEtwR3P9ToFP8tX/HeSnMuWVmExwVqvCMzgn0HsrAOoQv+kh3vml0oSGsV0qh
PDt8DnH7bhR7WI5oFLNVPDBT599P9z+06a7zYGD71SfaUiOhg4e5SK6p1vy2ESEH
u7R/wtIA6WHrMNmrmvJJQTT4xt2N+eb6j6VV4q3c4s+tx6arcqMkXSwGE9LCfwvk
MzhSod1SSeSCkXKhL3KffbarP4TTluccvgboBOT4c7EJl5dPU78+ztahxy4z/C/9
8uK7TkR9XrC4FSh9/S1+XPQAmct+FtgB23Z7MaaWoNAJYL1R2geIQ0Gq6remD5n3
6NooVUtSwycg1lnnIpk6WtLAhqZbxtrmlvV6H8hIQbel3lIGA9vSA/Ldb2WnRsPI
UzJ18VsETMvFAcoD0V7waCn5UtB7cmbxORzrdNytPLXDmGd/iVt4k0vzgz/Tj8Ux
Xy8Df+CvfXSEUA19iMJ73+VlrrD35lBWaU1j03dgY6NM6VZ8iZnK6g4A5Oj7Rv+3
KYP5LUmLUJ89OdkPoE2ftILtiSAdjN3xhRoWRKNeaIrQ6RhdQfAiF8dteBWvT7Tx
1xmo8fIdZ5tBgCVB9x/MqoGlOX0XGW+KCMdJpNB/AuPK1nd1TMOtUwpYdyVs9YOz
HVZhiEcnFpqHoIOPnsW16RxMbs/hp/yasYWhcjC69BeO0UAQEqLN9YmulbUggAqE
F04QsgnfCv8EhNGkSxFqtrtdV+iWVnoZOlcwiofN5IlYaxQPwvQxfL3DM+RxYXbM
rEwuu/Wps9BPrEP/ym3bFul/p3BpDEy0VZZW3hArQZyEE4lMRcYtf+jwT7Ew/JiR
6WdYDwEFRet4CO4/P/eenqoVr6UXZjaGw3/M8u+8aGiH/4Ex5tYYMPF17VTto4+4
dNwuUQXBe5tplomcSOzr4Qy1s4GMRlqFEoVvcrCeurvWsXH0Qs06fpTPw4U5/o0r
eJHbzt5XGiD29uWVQ0RP0MQnr0cBucuxYaQRhXTY6DjweY0Skb0ywNLYAp8sXEH/
IhlIkFKPr0lk15E+5VpnMw/iamWkB6Qj1sLl8dN3OCixSEsZkuULTZj7EaZq0PvX
RIDOIx1ivd7YUGMSM1GoNGQf+5upP2Sn7Y6pLI6CZmOYFqNeJMBrtjOM9y6QgnIK
jAFISAP3BgSKuocDh98HOMRUoyLX/D1WdqkMgt58Yt9a7wtR8kQljOm4HmJzM9rw
KW2cdn1z9gwr3DEc0366vUJyzs7K/Sh8aZ78CV3MnNtkiEonK9Tngk6Mo5iA8KYt
io28D6r6BoquuHARzDicwa+HwXHRO9/S+4CpcM714bq0wassg0SgE//RLZ0sNJ7F
Lbr5tNRCwYfx+8aeQJjqSoW/2uAdOaMV+HQw8aaYoNsrdP6uxnHzCKmvpQf/uFve
to04t/kdnte69ZlsTkgg3hXmqLC+qUcDea1bFUsLFg7Tzn69IiTxxKQBO8mWm/zH
Lnc+Apd+5ee8bXsUtb1OQC4Kzl8JuI61BOMxwiY8TrAPWJOdmgVbWPK6lRq92w/2
0QRCpdXeOjmBBMemRnLjKy7dyST0hogp0Pj59BCbG2YBh1bhHQ02tCc/rIR9xs/q
hFengvx5wu9LfjoTjddXpI1yQc/rLe2XsdkJzapZgetc8ezFjwrOwDoODd8z8+AP
wwp5UV/G8LoxHeIlwyS4SfZxWskbvBmWXfDUl7hFq/OgZvkd3NuHo8rz8T+JbXRK
2B3vd0FJ0bHEywTpxTNou6NWtsna8VbKTrr5jTIcVvEluCBpRArqLW/OrB+ZZzjX
DmlkKHkkJ/pmYT2QooQ4mW0rMwrAA/a+QE/HNPouhHbsKTIzj6uoLL1cRM33ZARo
0Z1aEmJEYMsji6tQecRv2rQZlVQ1sPfK7fuPzAL0ha+hQt9X3PG2BXwDbO+VVmGc
pTtCOPU2+zkbtl4lUDB9RE0YsFfz9eAa3UD8bWhREK0KKAOJ5nkYlDM7BWvoiqLY
cWbq0HJMGYgvztRPbkQHpP5ki93Kb0rQqevAwJbCFFDwp3Zaqb6f1WR0oYMHpUg7
SEH0LGCoHaC9vpx/mfVertoZ1papIDkU+/WVhsxkrhZ67ASxfih//dBf93zrFayc
KvA/xB74q+e1E0pgUPu1t85BZFeP/Jt8m51IAFO4pEwXhlPgrU34mvZB6osSqa/w
cOcc4i0AfwXj+mac8Jz39XOW1WH1nRUrBS77AX4aYVfZOORboc1xZ7rfIRtcpOJB
ix35HEpSLYUUv424NhPjy2DouItOIjJVZ7w9o0vL+aQCSyi8V4bSHM5aPkf5aomh
bCzZ22FKxcYOShrd1pcxvvUVUfWb/QhNr8kOyEVNOlGjYIbwsolwsb0PNOlIH9QX
7JUokDBZ9Yx8cYfOyacspXWu/44dhM1l8UB8PCZcp685fxO0QZmLfEBmZGwZqBbI
4zwFksNLt7J27Hv4nAc3HUVHdR5ShJGXZS0SLp/GgOI/zbLLauHMVb0rifE3NxvQ
qA2Ypj64k8LFO4bn9dUPzibBRkDSekkvpbiMlHZXOkFBy6bOTmGwnuJzn4Sktf2a
T6Z7LXZzor2j0jVf8COo1LAsU9K5wlA2CX3eyt814rJTdBeR6KaYvh9gC0FGhY3g
PlcrXvcpcycvIPAlfsImOApg/bva61h3bEKw574hv37ab6aBkhXcWgHLYCjPoHm3
GpemtFpjRYFMuCUrHO8y99M/yRm9QAScPwwFcDahzAoPw6NQxE5NEWcgCiXaZddX
OLt00e7IZQZ4q9n1sODRrSPaC8vywRqKs7DjtYHMffAFuHSE83ZnUlPove9Cv6z/
Y9UZTUjPs0Ac8TkMpfyoilN0qhGgMp7Q1xhU/5tE9LJeU7GDELLhDxRDzucGleSr
OMwxm9FClG+NNS4c0g04ppyz2flm85ZhbJr4lDrRIPmoPaMT1qld6EXVjs2Rdroz
NsFIF4aPyBjLuaoxC2do0rr3GariQODM+tKBawYDS5NRsmREP1iRStxak7rcZ44y
rhtGoAR0rgfP4GllNvKR/Q+AVKWYp4/kNvwptFUHvfG0V3VDHYJLNkQuBY/AUTJ8
Wi+VqwTQcuHnVnqkBt4ugQxcUxqk7XSzs+Af/og/boL5oKt4dBXq8dIqwDGw2ghy
XncHZsjpsE1ouKCKkzeCIDVXz0ALZLffaT8/DJu1fYps/uiQ6IjtS2ovgTuNTd4g
qMUMSiDnfDW3Ea6+haK5pZL5Qz4Vz1RQ6zxp+V8WI4dWWx5wlOKlgUdNBFHOytYS
r9YtIniCROFlWUVYsIMDNIoxIvlBek3k+A0V0eDCgaEG1aSmR031RKU+1qBlaAoJ
SPNszkaiowwH7IeU8M0Ie9/+Q9hxtXuxkrVQ/20kjliSH81i5/uLsvHXb5BofKbl
uGJFUP/3KaEuTMdK/5pflnWFTjKToMdBntMJMhPAokY8H+bzvv/F+2aZrjUSlDku
pcexq6da48UTX7bwVysphmUstY+K2Z+NbBdVunHNAmlyHJpjbYPWeFvn2wPmIeTQ
hnfhxYEnL1YRwx87WOSgLrVyqJDEYPpebHYqKg6hlDC+u+HEIdszb3M2XajvJbM/
VefTw6nZwCYtW47+Q79Zxy3zJj/n4X1XbULxDuiHiXrGyEMkdEaURcbDWzGsvY0R
NPunWik1tp1I+YBAkTqnH9KbJJGk48MiEbETIQSvSMH5BiXctTXRniNREiExd7US
pYBAlXdgOHLihKXU/YnUPGxI+a2RP7am9g2VomHCo5l2UaPSM0jUvYvhEa3PYMld
iuUURCqKkkATZ+GUjTw5tB155oN41/3ZdfFU8EKQfkuE2+t8+iYBADaaXzFnLhz7
IMxxODdVZutn5FsLIRBXsz0Y0e9HujocyeOlY/nEk9JU/9NARb3jwHFLbeV4iZrm
5lrqWi4o1O7KsY9f6TrVttDMlM7R7fllNfNARFRU6HPvcRUqbTsSoKer7aVjDcev
c4IL+ID4AGlIeUt2PJK8ppV73Y9tV6BBtqC5U9xVp4xSk1rQi6zxvQSxljFg1C8q
UJSF7/AYbinuucgiKKPcX60JnHM7H0scMbur3+dBOoRzbjqXOaLg8Fot3qMOG68S
zhNYCx4OZMgCY2YR8XDSqOcrekej+6RVTzEF6joIQe7vqSG78zA4dPcgcDYyIXXT
9hJSInwTzMeIOAE7Pnks/c+eGUF/fO96NLGi2tLpBBAeXZjGzFId3QF2wir9LxJL
wwcXKBkUousU5zqhi5GchSvIryz0p/DyCKWJit4iCb3P6B907/3nYVnfi4VC1yTO
eNPrbSAdDuvd4JtyRqdrGXWWfJQxdxgvgT1aXIuZK7IGlx6KZvHxHZN0iGKCiS+7
w8iCyzbCPkwSKAiEZOL2kJpYd257ULnKFtMM2r0H1xFyrCrZA7XqrxMhteewNKc+
O6ObGpn6CBmaXfCfHBQF/8KNY9ZGtQ/Kf2qm27CCNgsxDRPIvZhq/LkDhQZ1+720
RbqPPAVuCF1aFG9p6O5XY3pay7mLdE6dzxLpy/2f2rrpFy5Zkv5B1gfABgVGy4wT
2eo7c2Q2K4u0Qxh0iESvVgHxkERNGA/AUYDEn+gh+35TnH+lHTHzoWssYyHzPMjz
chxpXCN8dY4VRr+aQonvuXT4nsjdMMOYrT1LWv8SOla3hd9Y952gSEaqQ3pRZ9AZ
7ACn49a51bvpKeZj89Zbzkc9moc2EzKW5ALfARAIQ+dtMH1pfLEKUljx/IbGFwgg
wyX2eIsrpLdyJ9buYOrCQyXo3RTVjs8kA7hoTtMoi5ksNL9fo2pBrgTs9YekBzpT
28V9X93HPTHmnEz1txxTsK8mQwgLDpJKQcB5A+iC4Zn0jWDF0uGiHsJl9NvKMTzX
spzJmpEJ/MMCwt/l6E55rYgnNnfbHUyJv8BDaPgqOsbCBsJPqy1vLj8ZWFjEHwXe
MO/cFvaD4D6YMc4MTIsCxJbm8OWDEGtFabbgyyhxSRhf+Sg2erMOnAwIgjHMjVgc
EON+7QWS3fA4mdP5e3ZrOP0XJ6p8Y2dtVLhpXGP2EqjnJefvgOZ/5Rlbk24NixI2
yBZ9uJM7sx9V0PpYgbpwc9AewVRD7ClO3pHRbwH7C3WuXwpmzBus3szIC4dLKG0Y
eL/hNH8Wn3X8hZfYgyne4XDaepYWYO8ewtBKRGm6Bkgof40oddr5wXse7xRL1o70
1yed1eQE7skbDIw3RJ1aRCOKbhIe09yCQx4NGdzwQSWDt3knDhtD7H240WyOSOcR
cDBcO/o5z3dRKGOZYv2D2zUXJokWnauiJnAkLYDg+k7UB3cw1Qm9RyjG7ZlOUeGv
3eVW+vZ4Qu/N61zoHNU8TuNULBH9JIOFxrevLgdUAvMTWoQgAm0DRTaW8Uw2pNH4
UPRxZos6z3/k4S+pkq0f86g1k0238oehYLCRFfhVuSDxEOhHiWszbZ0nRAfLmeBm
ExElPOB0u1jE8GaZ9kHdiusrwxXB3T9v2oXQpH5PjU4J921X1oglGoDQ+GmkBnPn
1giLpiV7VQKKya2KzDj5WWYr+qRvwiAYPmEhXx/bV5jTaPHKwPdNHTU7G94jLJcD
ETCbn+LmLV43zkCsviA12B6Z1dB0+/oQ19lz2Xqt49RCI/qGRlotAWEyLimGK6kp
tqnGqu24rvhbMVz9HVo/ZNIeVh/bR04u4Rek83CFJX6Kn1iKR0NVS/zYhEi3JqqN
VjjWvo2j39Uqt8arQs5qeKMOhoRpu/GMv44BF/ajv0nBLhVdh5YN7BDZ/xp2WMt/
GQcTcOdQjV4a9BImmWKF4M5KhovKIdjK82SBEWmw7Z4G3mej0l3kvWAo2qO2oJLP
VIXjrHVFPIia1RFBi3mtHsk/Yqe9udgSmUM76kLbKo0xjvjFRy3OD1leU/IQ6Lpd
Ntqd0aNNBmOIfRVAYygniTp+SYhAhvXNw/bPhfQhWNLCw3x2mQdHzKUguixGtKEz
MI6eqNrPzaNED0EBc+JQGl34to7V7q7qvuy+g/lJZEbrArnInJ5q+ffbvYewueJY
AGRYbNtNp3nv2hTbcEJmKGDJtCnyUdq4vf75eKrhUag4nPWGEDNu2d9vWJdWlqmG
99z1a8EHP96t0JhiTLBrAMj5vp2TWyHPztdybGfRieCNy3tH6MhJFetbr9wijz/L
XkNT9i8TgYSMtFICRR2T30SY7aUz24is22R2LM5IbpptoxPClUMt2p+reCeNBwhB
NDy8rmTAJfi8NxaGn+kaT3g3FCHctvJuRdeJ4bum9s2pMPRbsYJvevWrIP/enFAB
R20/a4htbq72nSoqNsKWnYhmpOXXqDUUmypnmd4B7LSH6WlKTq89AYX0pGL7+zbs
2Yo1BHHe0BFVtPkKyc6iCabUBgn5v5WGcmhT0dX2MmMnhvIhj0tWGwJWZuMb26Ev
9t0OzAEJDnFcjTWdEoLu24tBWpkjYIGFJ5P6YDmnRodzEGC/DRVls31Nb1FZ7SkS
0B0Q2y9KMpnLMvDv9JBl4yYmZUiJ6TuC8QpEbf4kNP6cX63gDAtoRlEYl0YP5Tbk
TYHCfCJV2L0xzXDFRjpFHxpEeoOFdWvNjVEkuzfiRYffLo+dWLoHcIHfaXj9wRFj
soI+fbsSexZIm0a2fvO/nhCQUruVL0Q9cpB+ZplgwADJsYWLrH/ayxImRcDoxPzJ
T42SbvNoeeyMIZCfU1Dz3lYtYxPRicp57jCGASN5ZNGDybf1FymMQS5Yf1dj+kb/
VL1PAEdeaiEZfrXCARC2747qMMT3C89Y6YHdnOuNo7+98qoooiLNiXU2M8N0TQXJ
x2jqfRnURhkjoxPG6KEG8SMZF7kEfVl2Yofhb5mezNFx8/q/0RfNeqoclT0Cj/2g
lsyTdW1OF/9WaiVrcVUFJsIobnFdfcamQ9smnNmlQUvztZEc0Ji5PhSpeg2ElXy+
UViu8fNI/lRqhqHtHQ/aauP2S5YtKPQci3nL/F0p/qrvkxwe/RgFNtxvq7Gk77vx
rcktXVcPKURKwrnAk8azd4qI7JSfBicxI4DsqBxRvsUK028dViNKl/ocG/AuBrQb
83F6CONUtxSG/NWOHCwLDCOpv+8+ANe6slv2ZsW+zru+DfxQ8DqCt3kp5bErZU15
JR1Vu7IWHtQh5URvFHzfOiaUJAXZ5tZVR9zt+Wrlast57n8Kh8iNsZGPk4hGFCVW
iLS0dLcXmbhly/+VS1Z/bXiRm3iKMcL+Vl+wETzN9P0AAo+YLONExR1HugaqH5DD
iofOsK+ioBoH+25ihT+lgvrtHjEUX8jnPjDL4IYYLy0a2BAz8BjEAKYMffeq/s7G
+s1M/DiVpQ+wW1GQOYzshLWh9vhLVpf0EYamhJXeA557FCQjUve1HwuGHBpEAajX
8GlyRZ6TAcXmnfdzLCO749LM46J8fWGkQedarJ9IL3GqHXnJoozTNuS7HXs2mbpU
MrBmGzsHObGr2/PqFXb9+5uY9u7h6GKguhex3RL9e6AKoSgXzZCYL0df4OlKLEN3
XtTLmY0krcFS3Wj4ZKteOVJvxxxJfe9XlGwqPavI7ZesgBaqK5SQRDMJHF569nZS
+qemX5XguzmJ1ZWBfFBcSy4RBmfC/02epN+rNIlxeSeA04izKqpkTgdXEJHFqIHs
Pmng9tpofP2ywOygPMaJuqqQCCzltuwot4Jmbgud8/XV2IiZx9qwj1Q9y4vbUHwr
24bEY29BMvEK0qc5ofhOVXHKulU5lJdcTRXnDv/xdniOoG8f0dPWCZbccGJMd8ko
bzKcdl0R7Af9HoJzj9iJhS+8iE5UWOQmYiQ/E8L8ySrIh11GyxnZMyRNifzrZjWX
H64G8JlcPWmi6w6yr59PNR/9TGToT+C7iefKwfsgAED5uSuyYrIp3Hoz5plno/Uv
bCgVyho6nTFEU21+bv1llEvxFf7haOm3se1vMacGEP0WySYa8QnNAXSyxmuwmbr5
BVVaXjn23usIJnBB+Gxgz+Muk19OSIdLYkWSjlK7F8xCmebvpDtM+a1MonKBrOL0
WE+2LHlYq8HxfkWhMUmzrSGFSt1cK8SlcEdIulqWmfu83zYM4HVl+aCCd65mPdnv
NwAmsvXHXtlVxJLsMz7oPn6Vwj2SWlUkAZ4sN8elA3YOY+bhAAXC0XwbZgLPr2hY
8WW3rDB33QwfJzlctc/5JmKUJsHJmHm88CBSEtoM3yDyaFXxujFgRv1myF9gm8od
ynXo1zE7Xi5Q+mwBmK0e4G4HDQp8+ddVOfCCzlrHBiPVAgJgGplfRbQHk8t5BcSN
lJHFETBPJDLipo3oZY0bWkMdKGVSlTLpsI0jWTAa7vQLE5xfeQvE8IgZ6cgyLltp
pxXOCGFoREaJmY+7rZGOEP76Wl8BvEno5eIwv6rVyPhcB3Rw6XN5qJzAbtUCGuSQ
i0KISMK9MHZV3Ngohub8RZKIjWFpGfsFiLVjJt09/9Pi8Hgko2rEZmXL67awD57p
elUcwOURbMUKtcbzfQtjR3S8g1i89KFbZwmfZZZMhWydLqRfpW6BeeG/ru6rxCyp
h0chzkmIU/p/ehJ85Zo1Nar5GYkNzt3nsfaXN1e8Bu8H0babhbkZH7q4o8ZbvIsc
eVvJipE0O0P4h9KLsy/ZdQLcTLHGUYvEef/l784Oenpqx2LyMWFraPgzR3dT1//k
OsLctWoruRBNQE5UbHOfuttNdDCrjGQqDoPXLL+S7zVvtnF4A792OjtUqA4i2h5N
Ewkh9eN4IAkgx+4/KD4CR70+hgWGWHGd9f+knRRV8HLXa4IPkH75IVRU0/fTA34c
hJqaf6joQso/N5IC7Guoo96m0upCifXClT8nhEeaks+0w3V7h5M8Skit0YT0ynpJ
TYL27/NcSGaxnAnz5WBMHYheBLay99E5KPZoLGorrEeailaF/jrXy+qx+om1v5Vy
8nIRgJtYzTKkpPG/vtmhTkAnuEPDY21lM8gMz+UN069ZyG6EioFsrWVzc2TqnW4c
bcqVuZdufcBPA+MWdli2IQcmRgbHUDoaBP2zssSS87N+cbqWFzUXyj+ppIDbzZX0
FNrD7KOF7zVHueUhE04K3rbt7hUdTDbgNczkwlErHzg5DH+9GFvrnXOp08YZI++5
YcabKyK8siBPSDxBXRhrRP3KS1LEQY53Iiu4IKSgfiHbo8o4Vp4rONo7JzLvzz60
25FFLXC03r+F6HeVyBL5I8a0m28F5/0OrZFOU5rTr061oFw77o09ph9jn4Lc1rkp
irolVx+02sX2vmUbdOoqI8MsUPd89MQlLJ4M4VuhATAthNOiv8IlSxzChtbEwscy
ZFuQ4Og4NfHY/+TrrH17O+1qwHVixKROWne10wSe3dVJy1d1l5Z0fkiP3Yr45pdm
7uAGLfdWgFdASU5xpSUUf82dD0iw3JFtVMp+u4TdQkCGYhn+BAl3xwkiNlezzbU1
2CzCQJgdA94g045sU5At4gTUXT2BRYNMpNiLCvdpOw0WHX0dHkyOicBinnJYbqjF
s+LcrzqaruWsGCaJQHUBhmmmhGq5vnfvGTxyGzEn1tAgcG5HWDldPHTfqSdfIiuL
F50KI9UxOp/sh7hb6GrUr3CicGfrrFP2rDA0UpKNLNNB4pA5zqF2y7ui+OrznB36
tefTlAu5J6mwpxmV01tyMB0Uo/THV11vIQWfTcCfW7yfrI5jf0zT7DtJyrVhKKkh
VA6icRHfW9xUJq05V3iCdduXR4HR4N2B4IYR/nnypbQ31AriXb7exef6ErwBwHSb
xlBfDTV1YfKdmhzdGutq3KNLgXPajyIWIy38ZTFfENiJnCX7ywjWpMeBIBce2cSs
A2fViyEZpXe+nXHR6UimJDADhPp8YSNXzZ/r9iGUuJgqhlYWep7jV+BgaZeAQlRd
+mwmtciscA7v2Aa9o9bUKfKCr9NAhznAlzpf8Ch4bhCz8LhXl9PTFzxGBnqh1lvC
6xQ+gzGKbgKcfE8PY/iVJjG17VcPnKTxU+IYekAeDOUiDyYsRzERLpSEtPYan9ih
Cz2OKENbIKB9T/z7JSubgVps2qkggboDPUCDhJo2kUAk7ZQa3/UJAUGezebv5NUL
xjU8ZvTddUiNb/9Lfwbp9DoCNKDP+8HMOmac2QN73SE/G4gnPD6svARJgT03EcEK
EeVcR+OLe+fn1beXtDN2jOw9NMtEyaqMn65+FRq/0WPwtg+LcAG5VA6pdEVNICMD
tFFQQDl52ZDgNGTCnNRuVB17HcLQDy3kdZLrh0J87jyh3+Dcw33qD1jpuKjsF9gd
NomEoHyr8P+jApclwgjG0ugVcj1S1xSJCPTfxP2uMT9g5KRs39u9mwuSkdhlsCpf
jfw1Qde+g4Paxln9QrIHjPaJh4H0vfdvdiVvZW2MmehaZJjGU9mcCdEH9RLOYvvj
bFsXMiJC7yG49zPQE9cdlW3jC8t4N/NBnp84Th6Z8rZ3Au1Z8y3ajaknIPlw++II
Y1olNqxbp1nJ6ok6QF4Bnq42NHusam0KSFS3FP6dNZliIYk0/uHxIPnQltG46BFf
Q+0eAsRugZ0/InCUSZb5/WQhM1tONeir6kRmerlrYXh+9RL0AA6tzsVcbcuUoyvm
oi1722Kavs3embwONbgKkFv7+665b60thEvVrx0dWAWC2M/xq3ILxc0MFQzJvTap
c3jZDroOCIAIt3gt1ktx0jNQMLmfQwq6/CYKkLKNA5LhxFg0S1xac+odIZtaJzeJ
upp8f9uwmli/ItllCCrpR9eMFCbHsTcM8vuNcX0sUWzMFurYjxFG+el9zTcShibT
cScegzV0AANvzzE2jmQyipkEhhSmfrK30rzPZyQo11pkAvyFHEFzSVAvvGFR/djX
3Hq461Px0HuA9I3tVYAHv0ipImjXncHDLgyvJ5EadOy4DnNzhCdy3X+iIbTEx4qa
+fi2P+ImuyItTmw2P7+AH8IaBlEq9E/vHEm8HCB5Ql3QwCc/LmoExzh+Mv7mFUfE
Uh3gTfQw901K+mY49Q1OyqBWUzgIh/WTVGJDXYBIy40mc7mfN5rM+qeTN4+GEfs4
V7TbG3p5EoVyGpsQARH07n/RDdtxyLCaCI90ccyQ0OxQ6tmSz3/Bms0drKQJEvHX
x6fiZ5DoLl4lymKMFDkqqNE1K6480nXtL+GqrMFld5/lYDFoxfgYdNU07fRMAomz
varhr0M/QMqQEUuGo2gLwhtEFYhdd5TE9PsLlxPYQss43Kp8N5SAUhpVfxl/NsRZ
iOhP95GV4iVaVJzV7/YmGOVGCVHlwgZv4TM9c70hqT5NRXzwTDyfK4/CEtwl899f
ZwPHExu65hTAnvmHlwvI+Tt1HYQaT0aOji3cBNG+V822LYUYM4iQKgOEzV82cDJ2
IvOolqEhxl6ycw6SpeZjyqBOKSQIUNveIZO0NJHc5U1YrG2Aqgg59WJPQLKb00xD
lelRxOskiQ+zJUUa6amdhRJqY50luB9qI35B4MXjMcGx9AJTLWX4hmElfaH/CnKs
XGcr0hyC+6E3LtmtEyzlxDww/Az9fQqBklvV66BBDwnUyA4MhIG52ZD7Q3GLV4H2
LJRs+eRpyJ+igkTwD7XilgjEsjuh+T53LLbYLdmD5MdcATYrfwhElqt5Rd3f0Vgh
lXwDkukHqFa5JhH/jlCLYORJLnB8vi94Tu/mAyIYMzk4HrFMVp25Yt8mCLWdz3MD
+masdKK2Dd5caZGJJJ7ECLGuCut4QNq4PKqZX7ASe89pQY6NtHXkUZYcS22k4cxF
SoCtT0OXXum+oA16RcG2wnb10bl0zq71PjA31uBcDK/lt1h1RfmFEn9Ebj6ozkcM
3x1HXvUPg2YL+OOgv/RuFiqSH38t60Jl6yoRlzWgszxQ4WguqSLGJ9ByMr/P6QWY
jYUsY6J71EPAk8/9VkamW2UaB+I+ZdXpHTNfhlgTg5y7rxALi7NVfDig2fR2mdEO
9fyip9ldUiQkWcI4kx8IRWD5RYyBVRNxndUAD+TcU6wkorgDEX7x2TjG3QIvKLa5
J3C2gSrHejY2AtVPm/RhJmkQZCkw2Klsv6Ad926kSlQLSIOss9fPOIoG+OUhhoj6
kWhLfl81V5D8DNbuSaFpv/mElZ8HWGleE9JsQHKu5ZD+6irAWLW6lcYxGJkm+WaR
moE300tmI05TSazWA1y8qMO4QahdbTKnXPHj6jP2+qPpmmCz3kHqSfTL370ggDgS
Ow0uzUj8O3T8I1kta6+dCEtr37/F13AMa1OYGp8PH9xe5kb2rQjvWHg9XpbALHqu
DNeF40+DqyTyHWTjg1N/Hq8ENo+NYY2s3FeCvwKO8h0d2INrR3yAmr1ycRbPfWiO
ZHPgHdf+ldm7ezT0QL7cJMoc6CNapWVEBBeF8zvL++c4kDUiRA59XOF6SD035/Rn
WZvQd4nfTea27VanMJ9U2UE0X31CGx4qOQe8tqNvaWh+5rUT8zeKP9yeifdtvW2N
sw0rhxJ5FWzB1T/l7H/1u73RyAxXOsSXTQpH4P4THPyRk2RBhaO5Z7e8dnaGXUlL
Oixs7O4VRE0MSUXX/0NNAjL73tATVRc1QxL/n/wLbLcu7uI6Q7YwMMMzWnCgqne1
1UGfe+YTmEBioMFdNdhDbkjvBFouuHU4u5wYkvI85zNlhN4tslgKt7/gBusZXg92
RXKrirdDFGyurQDDI9XCo1i54zDKnJmwnS93tPYn49kZIS/HiQ+4bI1tHxF4hwid
nAyZI8Q7Lqj5KNCppXmaeYiZerRqK4VNN18WXKjeKE3qcMfmBq5+ZxN5pZTGkyis
9geU6xyn+o3rJ21rSkRxp/gPay2FyC0KKM+E7oFGTqynz4L7Td7F+OGG5CpUPMgJ
ekGOJMJPB2Ior3BtNv+yvLrz5ZQiAVWQRcz3wsGmJQWQv8WnHo3fYq2AlmgIv5Xz
WeK26dbWCQZm3ud/dham4GtGKHi+q7FsXF3Z8r57biee4ZyN03nARb2+LgxfneLD
D119USsGyPqNCDbfZ2DFoWIzKdmwnUhEV9KY1oR2zLb/jumMCNK1Rn/FzDJUctPB
kKCLweQez1hpKVKVXelI7Z+nJtwi9KWNnc1MAAXVyQNvR1b2bzHnr5v5IGqhPxhV
xoE/mjs4JSEDhF6pfi+Jly5RtlMKB+szZ7a8e7wedF1tkWYvNC/ZuVvJCytm4Is4
BLdBywCD+tKER/IA+rY8Rx6onGiABh6PrKI6OKVCmcWu8fhzTFYduXRrZxSmucIF
ZMeb9FEeCvM0MZkRTfNqtPrvwCuNtm+0Rf7rU3aGJihxbIcOYqDkgsbsRQmlEEH5
aM12oM9twkGF4P2LcwRXdax/hexoCX7odtTMu/KBAcCER6KxqT8FtBhvGtY7kyG5
PUB4ILt38nKf236AMmvskCf2tjbpmYLPmDAs9Z4f1X8h6aAfm0HsovYvMzAXirrE
IKrgnJ4vCKptRIysVEyFy06eUYrLItNK3M8DH9Lm//BfZooYCXO6ri5TfnyAWhUi
TRsSyQc0M2hzgW/BngDY4GRDOwUqBD48hYtQKE+cRnCSKBoGy2UBlw4zLEGIhPHW
F93+kn5BNK4NycQ9hi3iWNWf/nPFALCh1LB1G8aDeyd7EQmjdgGJPX1d0j8T+dTV
oMH13CiMC34Kz6Sas2Sc8/yF3PUnysaNERWKpvNv+XB4usOmjf4nm3sy9ZcP74HU
sQf46KjwyQHdLPeL0bHVKTDBsJR4lBFAkwhAfXPDB0x+GTbef0f1UhEsYiGR2ZwH
Ij1YxgHyx8zn0ao2GNTEsZPqKgoTko7clAhdqVYVS6Vdwkn+wkjALyi24yHf1Y5v
vvTgbNFomGTMrDHVkqs5ieG8k9j2+rkmyvj6gD0cXlbVw7wfY8AGxO7Qw2jXRUXi
3KfgCdeirAcrC2ZYU+bCrOg2O68I1b+bS5XVvlrwh/vtd/IHtoKwW/BCG2i6btDh
X3LXFobc67UkVB73HxA8nhmNMLQs+Mc1RFC31dE7cbj6Rxxj4DdjCiAdAgWABvOs
R/pg/Yl8pnjmitSlGRTpvUzrgpdaEnOq2yEHhHuFvtEKo5A0Uw2CgQWiHdCupzE2
x2jMmRKRcjizuqWFEa6/iwQpMcTw3Q7B9gu0SSOxxnOlB3AzGmX5wceWfvgVVWBq
Nu8cV+LPEtRh7jL0yhWtIUcIT1RZfulcTZm0cEo+rvveLDh89X8PyNmtBvPKGnUw
IO87ngzAOirsiTC3ZCOTzG2PeHHri0n9v5muU7qWprH7tZM9ut6kAVnkcnkJgA10
E0WQgVAcqllmCDl00iUoHZMXAUUreF1311T1A07jx4gYHuO+chj9W7FlS6mDbA73
YGdDXlb1i27wOKr5egKZpng4zwdv2kasB/pY5PtW5D9zjfIyA04zI5VbuORYvzV2
JJ0oS+DUGNAjPT5sAwbmHzOfQ0X5WtV3zZICueC3K4LCAGMhTiFtCaO3OMxXXj5I
CqWlIPLK9G5q1jTPqsO0ry7OqHFaBKsd3jkHa7aBzspYx9xn+1Sz9EDfHVIiSeED
LAxuBaWR5iyKNCOyKxMaFhr2dvCwSaZyRQIPypz9a8cY94JI+WvGxWS1uNQYPhkI
YzmfwtemJVrICXu1dNU40qz8EFDaFGQPU+wkAVb5g1jC4coaXZ4x98Py47k95+rc
xV8jG3WEQvzhicuv02n+jSy0SNCGAQkM0jR3ASsifS1yjxk2uFmb4np3ChMU3oWg
VzolybXCBynfDxTrD5nQEzpaE7Cmh+vowwUr/7yDoCPzoP+MjxsoWpN8e1+01N8G
0/bZTnOJL5fIE6EGCF2T+AHEwOouC9aK8l046rbAGdm2SuvPZlG5jXCRPfqZpseM
nPHLphS7809lPDROuWhTSptJZpotY+lnFnG4htUkJqJLGsrj9NMAst/bk1NFKfmw
c/89cGXrNX8sZWPdNOxHdZGssWWiz/YTVri0kETqw+6rtn43YloMNJfq0NDp+sVH
HdYPhfjW+WBYfaAdjv58no1lPRQ6560ucs227ucaWY8hXWsLYxAk3qfjNfmOFTHD
F+BBjpnvBdqehKxeXkDhAjui3YWojwZZmEPlkU0FdrGxzxKYRTGuRBjf1RChw6a6
QpCQK16sQ8LQiJD5vhNqMSsiQgKjgsLOPcR757R35X+83k2OajYyBuWStFVIea2d
SD0zQJJIR6xmJYMdEdhPHBqCwDmmuNskbjaVLp8aYJO4QCxoo/3s+uRKleJnDivh
wyfEp74JBmFlAeJSae2VFbYbUZZbCY5QWUl1P9syWcb0aaczUybS/XZ+31Vt1nT3
y3ijm3h+UPvkcl9uQr1tK2XB9nBhwOImFcL5ccXKnJI1XwzypbrKGZppVoIYDWbY
jgLIFGkzkXdpgAkK5xqlI0oasNeFIhBZaL52K3XkSMJQqwCsaegtXdpP3n5K2RjN
W3jNWaY0BJpQcYj2/4nwzbiALJbHwE77CFkGi67I/+zsOVLjOj35RucclVyVjk1K
jdAstFKfEihmqEpNflcuvMVaZiuN+1fBXeHksGNIXdDPj27BYqTLtDoSUgXev3sj
rutEIi5OJlsaiSabIJQH5WvpgvijFWsWGLnYtWbfBQL86ilXG5bVcyrs0E5Zy0J5
62m8oV4lQLL6R/3GcbqU6vlbysNFM1q1s0aPncUm2k19paabiKyC907Qa6BQLdN3
1HzM0KcpnI43G6wJe+bBsi1S/8vnVxY86xMsM0gDOH+qk4jUF/zjGqGz7RO1vhaj
qg1KCeKopMvSXKmj/AQdOw7jP559BKDz0gIGTGq3cFvjtl1p1T9JRByXaKY/icR1
Nwsp/fClDUD7tc2YuMi3QirtNB5JrQ+qnCIIWJIEgmLJO+Mn8va135WFq8I8U45C
7IR51TXsherC5Dg3Go1Pku1GZTLzlhaUuSlNPD6QHK2NMiEw3cRM/anLQ6M2BgDg
w8UJptPWvGFYNOAhjjcLJc8pW/mL+PMQWQzaolODEX0wVbFQBG+5hw54CZhu5lbP
SFqM3ZZThCe9yVkUhBeWxX82beKOhgJ9ACuBaFzKUfK2OienrGQvBK0rV3BIs/li
uHHctQDPxqjD/FweGGLaVGuLTaLa3sAebLeIV2a/cEjzkCY/zqyOBGDWB0vDSM+l
oMsEo1huAsvzawav9THQiqut/5OkBh8OT6+iChjT47ybZincrWCFndOhJa18uNO6
YJZmvkpvZPg6BCunupGU2Y6vspgJ+BH/UmxibaJyHsGHN3udkWTifoXGoi3c8p8s
xtsTU5Gd9TlnncGN2KiiJifOdOI6i462QacCL58keb4qBI7fDuRPOs+Pn5QDBn0Z
RCZunhodloIEpNSPCRJ1sNewtMPaLLRTKn0/HH4o6be29b24wsOTPKYEuanWJN5L
ezT8ZTHylUYp1dsFJcAo2ki5sYnl3Zq9YiHzGWE3HU4WHUTGrUB/sGCEyCMKzvjI
k7cGXULEXO6tOoX7ODilgPn6ZLHwxDuEF3zvXvRjS7hFzR4v49Y5/RgTV5CF32se
UvLjcYOsNSCSFhcC47s/bsY2sT2TOIgvkvoXOY8KDbj7CE5NTiKVZqIgwRxCy4rK
1Ktt5D3bNo+GWu9zkegDBveot3y7QonMlQzOLeVE6ZS9KMF69BJJnlRUeHbKGkgg
+7jyWHp1dCsiqmxIxT7xOekgjt5/m1kXthWNt6cBt42jvWiS2jktLXzQq/0atnXP
yJOxPfuutTXcC9qQrzhmjaKYcnOrRXUAyn8KmqmijNIFgGAI37B29onisqvd1CCj
LJhb5+Z4AllgDhsdG4RBC6RUpK1ZjVcL4Xo1haJLtOk7ZGZybHMaESv1WaBufvnI
CQc3rlaZUBGSocF5j0M+NxK6biB7oALGQPP2BP12xrdwFO7zT7H6TfrDGHrFYXhe
nsiWCJsdSiSGmC0DstjDCjMRjXPphHk6m3t+/mRKmH1UBzIsy/EpKFbFZZPUizM3
gsIm48YxHa+7oxjWwzP1WKpO+mTTWpPFBvJ/D1HKHU9jbz78z1YLSOA+W+se78HH
1Wb9tOA+AXVYZwSHEdTwrgnUCNOv6ndVywjNG1Lz1iP4jGt++8lY1LySTxPpgOD2
EwofW3wEq7V6+HQ7fIeX3zvQ0UBFjWV+JHxOgAIirv9VOqwtIrS+Sw3ITlG0JaoY
AC95HxVruefjhR1t1uR2PDt42f/qcnRmPG+qTlDN4FodFQ5hG2PIBDVwozZxa1EX
C7+pE9Fy6hLxiRBp9ycm7+B1gVc4ZqLzIv+vseclEBKJCgD1MQg9VPNc29ou1ykW
u4FFApZa90ly4CpcPII5QcHeZDNAWTGrOPNbTf5eTqrTlG28/QyOtW9zBMt1uBxw
mCiY+TmPOD9+Lyhzb8hsuBT2dJWi19sq4TKqw8LabfvHEJsIhEsyqv+hf9ZDpvDV
/P2/20vsZNac6lZis9q3z3Y1Vr4Xg/IJvTeEzogSebbLXAARtALj5EhBexsbdUMQ
4VKDWoOnbvImon0jkT6Mnhtvs0PqFQIlbT2YChSTSfgSr8xr7+t0KnGoRd1nFuii
mAoPFM/j9/e2ZRvDlJvwCC6JePmTrplMMzM4DnigmVqUtZ9xa+PEvVFR2rYSG6y4
I/vGu06JWNX6pbFGURlMzjh59tIO2Iktn7SlPQMF3VYoPAkBbq+rK85y3ghWTP09
YnLP4vyzIuyxrtvg1I1wJav4Xm4MR1XpbtZmJNhX31dnZmaqVWBBgD5iwK2Ss2Oe
Gz6Sd7r6DJ7Z77lbD6USoKJF5bctsvDNS3Vti4A7ij2s9eUWhrDy0bko7UbgvxS2
DOfrBsFt7hzfN7gQIw6gOWoHIn9I/6BOe4IUmVSJQ31/qKqX32e8I03Ke5OqVXSq
wM6LVgH8dBlpmVguDZr3MS5lk/aFI+AtGxu9nTNaTDJthfwyjRcH220IFUUTuYLE
mmNldudOw54huexGyVAGwRCTYDb3f6dHcaik4O8mONSGUC61k2oufCBSHC62wUU3
KgbP8n3McwdoXKTeO2TzPz3UJka8q2gQ3vgXY3PVLJoH+ldw71TsU8ldRfp/MWT8
D8hyvvykOIVTKm3oDl3qNQotxgzv7fjkslozeA3QT/BdbqZEdXO4uImMr28cccLX
kcq6XM/wtry03+iMpFZPNKEMHGaOlEYGNd5fpbJpZbEwpGQx1Yzatc/ZXvg+jT6p
dlmgSAbjTL1kpTVmrk7DIxxrV6KQ2q36YBmnQzZ4h4l6QMBKkkeywb5HxxDSU8Jb
y0MW7ES5sYvdJVynyWvd/B2X27t/85g244EGCw1P3I7KB2UZ4Qsi+HwkuHer7DGu
DKtJ8fe1cmX/JIGLPIEXiMaz3aedRB+5h6N0NW+tpvOB97MqzTFTu7zEcsHdHkrN
JIsjpGQyK6xmltnUKeAaQczcVhOE15lA4jL2bU3OOXS/kZc0r+p48bkp/Gy/LpAN
ElVLvFfRIwt7xvr7m1BR0kPvS/umJisBHT0aSNq0jwuKZcYXKBRzlDolWbV23sUH
K2WrFehcANXBOCziJfWdin4XhgGBIvdWLzF1udTwlTAKQ1Ftk/82UjwZYT3EcY7z
Zm13b1LkibKBQEOpr7UC4qIjkpU8XUXTkps8OMrCugkJ+V9L8c+Amm8jw1UE+csU
Waw4W9VtwBe/8+HFtIFWDErZ6UqfKEPHo1ogAPnCJgiLvzgPyrMPKaZ7CcSfpbmU
5ESi0ZD9sHrHIOycCckC8xeeH2KZjQRVW26yru3ooIvZ6qY8SvinupaZ7gjdbbK4
ON3xxKenfV2SsflOvVsL3BIDMX2KzjU4hH8chek7W/YzZ4a8uqIIPA5Cq1dm7XZh
o5a8d/sNvOOr+t5TRcPFBkR/Ew17mGdwFj9NfR2W1bBcLlaG4HkPunHPrFTDcuHH
T4xoWlZJjb4eHYuVxUvAFRi2Pi0Yp431D/h+5m0TnsIL/2rJPfVWQ1en4nVxaN7g
8tLdijLkL0hAYUS0vI5rItFo9ZAfWvaq81I/d557LA0Ss5szTYl8Wb2zW55hkwER
RI1pDAMBbyw9VM2LS/9SM9alr4OuJu8J0Ob+bSGqM0qcNraUddU+CPVXF/LNAcsM
kIZRHNNaihvsnX7b2kwsVitio+UnZtkhNZxPnxwed05K3fPeo559Cg4j6oQRdl4W
997TLKLJ9usM84tbCQULY2JNvRFUXs9rJZ4ZuwsdzOTq/TTWVXaes5H4fLoAUAwi
kq2AX46JZrQ8jXFmJwsIiD8KtFsoNKsekuwc3BfotXaRYGkicVKBhFe4qPBftHWw
Y+2FJrVeT4PO1GczXZebH0Dd8vS9TIZwCDaqFWe4Hag88gSCXmEf07c7Wmchn/Zh
7WpzvVnq17sFfixKKsD1j8VweAZskbaj+9e6CgatJmnrBdXgcxyLLLvD7l1MjmRH
OpSEzKXTirJs3kJdaY3eg5wHWOxxvcm9M4LrRy7tSF3S6SYhIWSdAfQtStPD2ZJH
YrDpupAtJXKZbEvRITwUukNKiVs3hME/gtOYjO8dzscU/s+tmi20EYsSNnfHJ9ly
g1c1tzJ1V3tRd7vzvDd7g40YLINehr/S1p3FvFjUv/yWrpmcmUKHI8Qku3hYkL0A
68xh7kse4Dp2AzSm3Z270lTX/B/mWD5+hKSs4XK7LtiELQBztXEL1RZUCX1u2CSV
OFkLpjbQlym+kaTSyqz942khhwGbYyLOqsG0oYqaWy45uGDJ20KaxDlX0fwL96aK
bn8wzVyWqXanTW9ptjxZP2LyVSNWi9blaQzfZ6JamiIoWzdIddWoPOE7OxYcK2q1
ZxyES/EkLl41uayUVoKb9/N23LJ0cE38ByPqNXYGxxUBuM8y76eZ23KJjFMMir+K
+cVHJRstTtdkjGQjU29ZDwYNEmzyq1xjIVsKK/gMdwbeG//Bb/EglEymrCwaHOfu
i2/pzNPsQamd3NFsYJ0cA72Jbu/WjQh/yuY4RBqDKxu6LtQ5Zx+rWBj4TAAOK0bW
Lf2xCbUONmuyno186+hb2fueaHn8S1wJ+q5RHPxM74U/+4i7DFm1E7yZzqZgzK6D
r4k/OBzhzboUDa1RuT2eLzqme/j9yU4GbfG5VMI6KFj0tlBDM3GPa4BFIa4G3Iiw
jsybNbSgmfXnSbiNRKYpfU7/ib8ucWZMT+Nh6ngBEFhcwFnDgncSAwNS/3BcY0Mn
3wAzDIkb2NXJreTA1aO+in0r81DATVkMRJxpN+0g9Bp6w88q7Tl1cIETWrQ4pjMZ
GNArDmbtUbCdGAaNxIcsP1P99JQJdYuk/jWxvzhrRwMOxAf6LJTprcFNypsY57Gr
lkupSAjFmFaSn4KFazutwfaQZ3dl2KVIFbqCNN6aDBT6QafH5uS3DIG7Kb6JkJJP
csd0kj1zuvlF2azqKkd44UjN+LUoOsnCQ2aQVdJguxBcbHk26/H7u4fRNzM1Y+zD
QpU2aE7QeskWVnOeUN6iOczZ4NIRzAzskFUXDUu52E83b7hzMGJZh5qrOs6JEK+z
2y8DKv+QgGnzpgZ7FFF/R39JOzlrwfv9Q/KWe/I4aBjuHoWElDVF7OBkNipkWnAv
r7oe7Kbo851hMHs8Lli9Qv1lWF8u0Pf9z8L7guRI8S2SzIjge53CaoTEixaZkpYY
fnsYTsiLNoDypztY86AXa/irKk79xTWIa4rt/KMg0ijgEAwgEK4T0SfvBfguFyB2
q7r+zMu47N2WF598As9CaQFq7hF2aoSZHLpfDA7P2yHCtLMLdzDS79P0j0bbIr0s
pI3JxeOQLy3lGzxikoT3hv1fTP7HOiL26Mc6Y+AQrsL9rrR0seTv6VfbvlWmngkh
QMnk2Yx/r2UlUfcK5eQGNPtjYqrFtZlzB0ITfMl3NdptVFkPEr86BrKEyja1Ae90
N355rSwLL8v5zVJiAzNzeJD8oVChr0DvZSdNDTA1nlmBURjgmmKn1kMEGP7BJ4+V
LO63REuWmIfujhCPlqjk0xX1JpfwpMYUNGbS4AYgQMYOAOM7lUboeaLf06UEZEVZ
NbF7eFsd8xk8WgoIuKuEPxtCyWFPGzY6oGTDOuD1aboJleG2z0bnGQ8M4cM9/nNO
2sH3LsFlgnIJ/vik3D645t17dQY4vRpVBJBWHTX9zHnTk4xcFgSHes3PpsuwGbLy
nQpRCPb1x0LEQCX+MHl1SiXK1bwBoEM3gt6pBLUyhnbTCRFRhXQsFavxm9kKPWBU
219ZXDCmpxg8V3BCqE+g3V6uRIBIpM333aNnMuN8UAIHtoxTwfqos6t67BkYweyl
9UUnxopEeQJ/4IhTfs0b12zb0BWT+b5HdiNd+OugGgqCXR+4WKUfslkBCdEM41nd
OD2FdVxhlXfKsO5Eqo+QX0jywOOBujzUsiteGncFhV4YKlO+dBHrBNjKQUfsKUFA
Ad5x14mSfnsdtmS6mLWtW/haG/I4rN06Kd2LA8O/qv+GrqIH+oPHsqLeHDn3Ntm9
MNV6/3zfMiRel7M3m4bc4ha6mXoB8zytJ03RwvXgv1oEu6XNyJYggO2JizsMziLV
ub9EEwxGmdFa4CG58iF8UaK5F62tPf32fbbQ/ccnh/eHZKbecLZGLdU5GqNb4kTt
MSxdbs2XzyShGWNmSBZcar1gz35N2EHYZFdIW779G+Nmo5pFBsVlnniwRSNi3J15
FP4AsjTfRNl58uHBSKUtJxfl59UhTI6xxTDYWDIiHFXTjI3y5NctkRSMfCYexF3U
CJUNXK33jlowu1Gmr3RbJXyixqhFHi2mmYTwBG7LJaTU0CqtdYTf2CfHKYrD7Rje
mDCemwm9Mobcc9/ebQfCJZJwvOlkWuRiCcBGdhTWUGuGLtWSkIOVEQgOC0y0Dwwx
1Qs0t7nlE2H2l2ZNmvsDemWrsyTHjczCHD9NxmX2NOm4CglP8XFfN9/mBd/2CmJu
kzoPDnX8053PtQT5GQOsxgqEJUBXfv4OZR2sMePbG5PVO7uJcIQnZ3HT4tb+lvIs
nKJd8UGMBHsm4DGbHPzqXXKgzxNDChxWh+1YCx5hW99rasPGzxvAvyY1kGgjlkKJ
FHr3LV0MBU8r/4NVaNBnMV3e+J3OFW4ZrF/04T7Udjk98MEFxnsizrfwRjcNMzNW
BYFpZ62kLazkbETcnpTGd+M2s7H6iTjVtPzL3klgthxtjNQlUv/myDSo481F0TPK
cDd8V/Ff27X2rje5F4mnLklFdH+KDyoi04oPKP+yqvYPo/gIdLlf2B48H5XzxJ8b
mMWYjbLJZD0VYwxMoqDa7eaJUH5Av30jV1zoBM5huG9lJscNf+H4Qyn9za+10cMB
lL5nxdcSrbzGzIEkLforISXlfbmP3gSCihYqsopzpK1zJKNa+H/G8665EgB6g7B6
qmRiZYqREg0z4sMtm8MctHKIbqd9vEfK0ylvtfnFg9cVQNMT7Vi6FHqkNKsgBiSX
JjRRlv+DmPmIdj7SrNIgDw/plrefoMaJSOOdNTKonaqLvFAdzGrZTGETtB9oc795
UKqhcNLcr2Yf66nQDnnxTCgNspRlNMzzEXM4pmnmWlcss4xyrWvsdu+Kp75hD7eX
gPGiY4KfdKnJwMOmNrKf1pYmLN3I0TdMUNrjMu+WbxLFYKS7ZDlqAAlWHu24zJdO
0U57v+qONrbZIH/FOCW+AJ4NDgi4qRiSS/vHIIqUVgLfprmOKb7oHqit7Vuly9cY
NV6TkpemOAsBeDUFrvN4OdLbVxSJr86NQZDa/jkdMb1YR17PUx95stlCEPBca9O3
9NDQXKCsGxPp10YEEuszLJv1UKQwhSFjKWDHru7bR5QlHmOB196QiYEzzOa8a16F
KQdjJRHT704Fi5UKANDPKCnczER3kpH6SI+lt3rucMrAOHcz8IRrJ3ejIgf9Ga6n
eIZjgLKWiS2Mi8fe+HCrI7e7q2PszYC/tSrVhI1caMEbHzMaQFh9nzHCAFj6QjRo
zuT7ybjMj299tO58WeKY3yDucpD0xzV4nBi8vGzR8IrcJmcU30BoaOicUrinBUS9
lZyTUIeoPE5Ldpbc7YT5jK7dy1iIo2euJ3pcRQG8s3nnfOmbvChwhALWgO8HHxe2
uGlW6Fd1ZEpF3df3VZcMZZhtKl3cFxzpSYWk/BMH5qczAOF6nPCroWJ47ES7jg56
745A4GPRJQSMrXmAZa+ESyQL/QiAK6wjRfT7kBVI3KMe31X2RNuXT3cYIVowOrtK
uWA5ITpAa2k2lIABxZLjcQXxJNGfWZv5Q7A/ODzDqmtSWOeOJXTdHHgp2irsqBez
V9gHPUFmlBW1D+hvWs+OzNq3F3z7acxFumuFNVL4ppdQNFbe1OD9UcsVs/M0C9WM
3qsESajYE/XG3xBuNaKb1DSbTvWlkUXz6XCXJpj1CnTiKaiX2xQv5VN0Yt7nFSA6
wg94DXJQ3Vz+3qIxlfLscKRVn3swFh736YAid0ffqb8MJZVGCSQIez83xRL1+USv
JGa8zHygIjRQzA6oqKvUCOVQcXnGAuPLIOqEGXH50A8Sx5Pxy1Ya69qxiMwdF3QI
85//Q0AT0wByF1nc7zV/6oDLscazWn0Tj4h8V/7n7CM77gTXy2N9MNtjHycqaPvG
slfV7yOC/JQD6/lY6Bi9uuWLX3QEtU2iBlHoO3uqa1CZvfDoiKkODCd2C4YTqWwh
rsFMVEHMPK3zPbKnKMWl/DaRvmUo906eHAxNN+A9leLreERfnKY0vW8oaqRN5NdC
TeAE+Dc+gjzUb8tGOpHSccjN5dvgZDo+tYu53BOIu211e/p7nIC2wEVNefk4BD4N
Dh57qJZ+iy1pE42NxIigLAQreAa/9mbG30PzL7QRi140Eg2H2Qe4YbH14QoaztMr
zgCq7O4dKdWcTIaZTCHnQXIlDTrh4AXqv3ylyps9YcAnO0Lz49u8kIgdE7226zrM
NpP6VhKYqrPF/eZVQ2XPWp0+gMji35flx8MhqhNtoHCWJOGb78to72j3LSP6gpic
Ma4O9DYtIq91RdMdkPs1kipH3FnDbs3Ctl8gRAEq76m0aExKAID1RHRfPPzvifS1
XvN704qo8Xj6YSlxq5kTt8WMrgBzbDfUyme/UG00tfBwiEltgY6ZpP19tcKSZRAb
XvpoTi0CUjPiQ1NjDXxatbg/tYIUe7a1ObvG0v23HNemYHUgmaa11B1k0vfHqjYl
bN091Fm2+cs7ugxXpSR0oHby6lxwJ1vogXiZPN2mUzrI4+CBKWH3/Kz4jsrvchMo
oSVj3OXXvYlQyDKSVCprvzc6spKhk+lppqbY7rj2+HDbqbvms1PfeByESYT6PxWk
UD8Jgo18brPD76loKNuRnFDO1QPCf1i+yxncsIlkDk4cxTKA++hb5u7VtMz5HBL8
Yos0qai2+k6ps5PfjpOTYFqYnpjhCVJlVarXl0f8RTErqhBmRxglEpSxRqqQ4/KY
sXT+f+gMfeibicDzRiHV1nuvHkzih+mVuXQfdM29Rv36npqeZoT6EHfJTLM2M5OJ
n04zOqQZfVaBZVeIUhto7l3VX+P8XzcOVaGmR9P8WGlx77c++X0vsAdEpQGS1MC1
mgPMwVo2zahOudJC8hxpgjbFbH2RhVOMGF5f1yU/6rtSYY0xn3H6xxmuuuw3INNd
4F4kZJTjw1TDNXaGvl1y+pblOxA6ngXLQfbXZeo424WHZosFqLDb1Rm4GTQ59OX2
TX4qYexWHFmsJZWJkpZRghY714UlmC2CJS4kywqZNgLo/NjxSKZbeQhAfmYXWhb+
rtrUVis0y8OuH529ww58uS5zEH27miK/eQESsppNnB+6iwGwSGCLANFhiiFK1M+X
d3Zx9w2I+BUvTr3eoUPAYzzsMSJoGQ2QXtdFLq3HzTHsDdpLmYpjWafSKHTEBA7B
e0TH57j5F8ytcy74fWzKkKrKBNeRa7GH4XMDb+Fle176wXEEntzPBSzvFAAFHzbN
e/sj4aqhL3jyljdZWD+p+SgUTYrQ4/E/mXBuhQwLFVKi1hBE8UWmiNtHgcDMfKVs
IACjLNsPKvsmg5rWt9pW9JYH3A9E9MlxXIOaKvQAhgIyhuyusL8DudWH8/CB4TZF
QRhn/TnoZxtbJ4rx5DvC2TXjrqR+4KGlx4liWGTUHG/kR0FWqO8PXw9ggW9RLEaz
WtBkKxBtN35lcq0YDcZFAtEzgIYtSrPFIrHo6qGX9eXrQjwPZXVouMnmZiRiqg11
NJegV04fpiIMT9AmU7wTO+slrr7ry5TrAUpqSu58XA8ml6yUXR1C0Hj/5P0OBJYQ
brbY9QF4mwOALKZ+qZuoGK3JVV62QiaeR3g6RvVgPBHF+WzyLtlt1qvibbU/8Fbp
5xNb2qHbcN9ymIxAr8uvaW1HJ2rFdxml805K3HHkSty0bqL3UGetIhnJM1Mfg6Yb
YDMPPUqTdrG5VJjn3/rk7WiLj0q6E3jbZ1Zd1pFl4gkAnPVJ96kye4FnkvZUMVV9
2x9noLYzjfE/mYXZvq7K0WUc9urz9/9S03QfIoydO8guSn8b1J6EBGYkqZHAyrxQ
oszv2PBD5m48unkpIJC0fgCbmpPO7oO4aD0To3vWGuLUTYRSXCJvBauInLU8B9rs
FiZ5n52wgHsBocwciXZNwoz1HehU1JjiBY1zRRiujShM6duZEyN4UqjqTu6nUAnH
Bs5/lM5xjhYTsHox+unsfmkl6Cpw8OpTeiaJRNo5nylNX8spSYBg6e7TP4RwEONj
qlA1+BKFHSuEobSmVVFpeIN99ghdVTWa4OAcdgqRtrKNa+mvnsLbY5Lz3p7o2nw6
zB/wL2HRJJnA/Z5K/GlFHTP3Vasvn5aenwad7+3DwWlMMbiQM/8lYdyHYtJd/GdN
TWRv/UP7HdII0gHPZGLOJYsI7qXHWbSlVjcLSvsBEJD0TrcdwHZiHtvPU2vJg7Vk
pMoS09mJX1GwdqJBvsK8LH/MAjhErITzLPA1AuDfJ1+gbswDRXDHf7EJV9oe9Igw
av4cz20ZYjr50pZ+eFe2++gjh2Xi6HTQ3BN17vQPZNHzgfh4pLoAL4OBdSftWylt
gxo5ouJLfGsDr+2gvoX1Q/vNgwXy9p4RLura9GJEdYGl5BnHVSiKVkdFz0YqMTdQ
c0F8avvLq1ukT6/tXQz44hhIIMPEFvSYhmKHfjqcPijPPqcrvZGr8BlBFxi6CXtu
fZ+NYYgacDQUr3UUQODh/GRBfNXOPfL/A6CiBJzL05Oj8D5F40jr0tbHvu7DljOb
EE2Vps18FSTlweB+jDNplZm2Bj4QCKOfrzXPX1awEc5pl5F1tqA9VAit4c/HFvE8
uOEesK4GheoOXUhDjfqJ3JxrzC2OF97+KQrOGh12g6TNIZJmKTNtDGh2O2oLS2Xx
MZSFg5/JievykbROCeS7UuU+0vMVWKi40UmOW47w+V+jQ3a0kQKuZZOQQmkTPCi9
39Cv5T8MF5mw6ve9EzFbZjZTrLInR/WjxiK7xWObv9/sOPRS4m6BBVTmqMvVHjwn
zIt2ee2SArGhNBshBImCOklLTTvGfILjTm1chwLhpIgK8NaBrCVaFH7WkIUn4yx/
pm4E14N5x4+S/3IgBboa/284D78LfJK22s5NlKdTvMISe8nf+qMl45HYYSsVgwla
03u9olicOnt+nCNkKNBsld9PR1bYeyZDnBqihL6g4OiYyHG/0AIiMeRG4S4BRWuP
xsNL0/b6/XH8pkXWKqYyJYL7gpwoN1o29aWH27Gq78g4W8E2M23Nqwf3aETvn+/2
ySx5iHEbtcC7f3hF26z9GcOUbLjdcvu82NG6Ng543sFGL5cW57H96G0DuHIofI0a
/ZSZVxx3gV74nPfwL/TbiL7UsI5A+Z39VHZ4rPqHfI0GFYISLadravkWVQiphShP
ZJJ5Vt4hTF6R/rrjbs+PH9biEizrnDP0fra6gW//Wr7lqv3I11ptgPQCPakt+1g4
Fxkw0qriR5sPh91xZz/88JO6M2CimTAnJT0XS2aIxUTnvbm3oXvzPhW8wknhZHze
+AN6g44NA6jvtJ6cHqiapMqzZM29dTlNkj+B4eJVoJ5ILVbfyakKbvzu1hFqTHbG
7VDiaLi1Z9KmW3j+Q8BtwIqqEITFFXdTGcslLNKkU3EkI2d+juHU/Zd7EmYeUgSs
eUTnAQtstaxtcwKQK1oyqLNdpI+Ry0JpA5K//rxVaYiuwv6gs4lA3BNdjbB0t9e6
ec4ywoADacbO96pWN2W1Puz75sGoLaYNkMGkyDqVgTzqbdrwlRaxJDz/HUVroe+b
aILMYAUte9WsWzKe6xvZF465HWLiZNuBoAj45quwtNqvfwho/sWaxfAUNLZu2MzE
pjCjzMBYB2+j2UNO8hlNZPfAqmIaDY5YX8/jTa6iPMofw0Vw89+F1EIc4R2Zes4n
P36XaPm8irBocbeuukclcX3b3ePGg9BzUCPrFJ9dWd8aamUBwGMCCnZH6OSHNFVj
mBNYD9FdNxAg20ODsx8y6zF6NdzpwpEgk3BEC92bSpckp3t03I+Cr3BOzaEbxvAv
9iSZ6ybK7NzNY+1YMWcV1uZXszgWiGlSv1pTqGj5lgmdODscXDXkGe/ThNOXWKMI
Z1wfMVVdYoUrtBu0Rdmv/M+tag1vokMNgoeu3wsrQqMBbi1j5BmwLXiKq5oxYXoa
+amfhq6CXNdxSSgwhKzGc4XtXF+m1gO+1GJn4kM+wVJY1cdvMBUYH/KnoEGnX7UT
ZGkEIj+yFfd9Sw4QnkKsYY2EdflM73L+Ae5uwOUB1oXZ3A+0nSSsjmDQUahs8ydv
0iNAkDSZRvdSnRnoOFU9C4uFLdx35qCzyToV986sYx67gE3s9GDpr6ytjATfMsEj
k8hFCBPhzmWexhRsTsaGUP3lrYosjsGfqQqEz91juNZRQcSc5swJS3jni3pl1K2F
7HqqlkCzpYWt3dn5+Bf8yEEcE/6Xj0PKVAp+qRTbt18CDQhaPBaObX04wus18q3x
fDwEkLxEQISyYFyqEW6S93Qhyr5K8lmTCjuytNVws5LR8yDg3t0FA7aXtc7DP/Zr
3SdTZOkkxg4DmPtZLZpX/Y8EWso2vQZEbatXkFU7s2nbXktvvyipoveg3KhjxyiF
ybEBTyduM+piM2YsRZxVPrOAiNMNDLS7WpspE+3IJaKoIh6ob2ts7aCLXMCx8hOT
OxzFe1yIn4XD9BfUuQV6W2+No67yBKNp75WfN7WikVs3KLeI0gSPo1bE99NSXGGu
LxleSlauB2W8LuShBpTCufKnkWobjVvQg1QgA7+Q/jtFxV5z+splLpTqMhbzhte6
XJBhaaDlXnPVa0ZrX+ReXXCN6Q7nDpgsNjrUkPZHlwBvdSnCjGxu1W5zUwKQcMOc
qWRswQR9nEMUGqEzHIVY99cxji5kT4pu2NB69z4jJtZ0z+6l8UzUydWK3LECIigX
JphZjXFWBs1GbTsmdHA9kQL2K7NP+AwAZlfs8y9Lcqyq3SmV8AWtQe04E2M90TEl
C5kQaIYzzcKwkuQBI+uSNxmwJRrmc5lNPI/W3iDK/uWELzfT6F2Fa7Tm/DTw3IN4
iE8VgQQ+URZhkunwUzjWQ+aqa1s8fUGft3nGtdUUPBTGYnHCtBfHhJyb9KSiGcKM
F6EP96vQu9n8+0Sit8dtFnbztov443IdpsiR6cV6+Xh/+N5bveRox6UJ0/vSVbu0
7oNwDSzut85ZVQaI3nApSOO/bX6jLaUwnrjDmWiT/SVEAb8YnFaMvDB2K3mLGYOR
DSEJWvVgnZRLwmi9sqjTugKj0gx27Gl5tm1Xa+diV1GYSDpEz6boHuWKhm+2qT9+
lubYONMtMRVC3/fTTuObGb3W0OIg3mD2a9FDbycbQiYZedD3zM+rPeSG9q2wfjjI
ZpzxYilau5F9s8ojCLBl8+NMFMPmrsdulWDo9qJnUNg0SBTHsQuPijSOn8Ze5mBJ
2CdrJ2piE/ekqiLLS+x9lLmrwGR08EaA/oUbF7X2sjrSaPxtxc9Um0uCra5gZFmT
9n9nmgDuaF13ti56C3YORzA9hrxDqDkntqzRBwKQ8XidkY8Dawed2NnLHh0psw61
Xanp3GnaP+2uQ6IB/EmAyVLEnO+7Jir8uhwlPP8evz1TpefupRmER6ICQC4jJxFx
zriDLAgWR3RGxW08yfj5NuOjelWU7lHoQmvc9t6fiqbYS69zdFhuVosTvMfBNZzp
V9J7fzneOFT0KyMqtu3HoR3KGnH2co/jfVXguGIgG3owKM4vc+lfMUua4ONekwWd
1SBOn6Hw/mt02f39tDcVMV0+o1zJN1RplK+wJSKAYHB5ZmznxzwFvFHOu8ac44AU
PPCMreT1MbRVOd94hj1Fmum9ktQWoChw6xGHi1RQqRkyJfryPCHT07yGQb219d4R
6uGq2ou46PLHIFEfNOZIeZSGIAZzCeIobxqWxDMI72uX68R99fj+wtbkomUfUHjk
w6Vz967383BQwBctYbANGjbq2vhfu/Zg9qxMBGZcGWiRhnfZ3SefVYH2z43UXbvW
+fH9TdN/DNcg/JIEvAX5r0UkJc0gu2japeJMNYXs2jTpFRf5gCukgmAkb/f5NbDI
0HrDjc3w5yn6KXjr16OIl6JGy+R2ELFmcisWHG80Vnp98kAsTe2MY7vQ/E+FVCFI
VFJv3gLCfDfsNNd+/HWX9oQcm+rBYscuN3UK2FFrufB7uudrZqP27FFxDFx2knQZ
wCR5O7j67/Vc/rEOgifekzxWRpE+lkoqkkURqM0VR1JOHNBiCzZyIOTdGV2Tncu2
DKw5MT1NfhappfwophDc8sUnd4Iq6paWl7O4LuFio6ONYbS+SNgoGWvxGnhEoBFR
n2eR9qI+O/F50jr8JHT5UUPHzC7MCdvEsxlDV4JYOyBb9MzhrY3BTYclNQzLU2Cq
Yv1PcIVcs25A9/tywnPEl9P8v3JGncd6igYkRi93CC0SHQOKVgsNvKwVdYJ7dEjm
5xlFb8eRW0tfMBZQ8oitnoTRshA4Pxj4e7tuOcEQLkqzqSzbsX2+kC+FllFHFQOO
gqMC+fnSXs/oMeBbmuI1IPaumMGF2sCir9xYyXd+WHDVN8jqloJOhL7iYa26ooOE
CUImTGEH3ou4z+H4Uc6wgeGfb8EOQi8fnSuZUrXMcJgzKcXcEhU/k2ae8NpglwTD
8arrGVRlNoLycKUJqNal/j6bSarAXpQ9SHZLvkPolKOfBKTlRd8GiuTl/TkraWu2
eqRipbBFOKz6mqV/HxPNITcNhYxyJbAcwzLtl+WXt62JeT2X1g8F7K0SVnDP+VN9
q2jxSeaTE1wJlbpP27aVv4mYYV9YtW2HN5zEdziHW7t2mv5/yJK/twe6UF9Yp2aw
JgGf3sfDhcA46FxIpiQE2QKJy5JBA0rHlUM4wIDW+YITXIgrMrVGstOez9x2z8wf
lopvGRfi1D3yWoBFfp9JK6LJlypgZlveb5BZ4sKGN8tLjcL2x9vK2f67FgSufCqm
BoTn03Y9NMlVV5XRgKLmpsDtM+flzJIpUqfKvKzv8TNUglyV9j2TCcT6uhDdj2La
z8IIJX4Nyfep5RfHP5T17j7+C85f6MP7vOnjDu1+5k0=
`protect END_PROTECTED
