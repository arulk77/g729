`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLG3o/msZ7tVyteCbC/CYlryj2QZgznOJ4gIr5ovCevt
LNCEYGiqxG+INb+uqvRJg+O/eC8AEFbn2cYtYTXVF70D6yef32s+eeoBuscr+q+y
E5rcisE37m+rJzG0jlhLUXrSpqAAHctCBHYm8+rY23yQPLjRu2JPsoLcqNBqSXkL
xdB6QsZL3Qj+ljVzFg/FrLnPE7OD54RfTTw0gyA8Cp0ApqoA3lWi24pksPYbF99K
cIgAdLh+2YMgPT5maU/fa+DvT96wuZiJyd4qUR9gjZStU5NjwwmXDj8N9YjsCQOl
2mM4Ibg4jJNXY2JyuI9tmXN3IM0ycCLpy9Slr7e44IRvv9PZ1xgE6As9wDY3nUrr
GV9hgRftWkYuNChfogB3DTZeeuZ3FTyuwrbfVoYmzZEWxvdXGJmaZvQEADOY5HnX
IlIkYeyniCcGrnvkQWy38rOZKtFWjMTkx3+cyQIQMLQTybEWyfKqh04Ko5vOYnDO
be1LfsmD3Fj6vGUhTpjUjRMYaxbrJjzUeV52DsyrbIJrZ7/+NNSUwD8kaWRSaxSS
aIhOoeFiJgH/LTz/yxnBL1kRnf4aZP0DUV4LmaFUek4sIlwWVNJUxwwm7ZAFJRxg
y6BD1RPrMGUO0VSVIdEYE6tikvIn65Q8FrJ8dsIBPCw3XMgV02Pjk4seMsJPJT5D
XSvoKMMT0csLPBSXHeDbioaDgMQOC4K5yIaSGzal18f4c0kZERhuBQR7ZH+zNCJG
XkZcO+teSbpzR4CZx5Ua/7jwlK4EhO2m1yfzWl6+devhB5eckIO5svqEdkRNR0T7
QJ8ia+C+6P+bfLpABqoyBf1f9L3Clk2mLDTO/J1GbKI=
`protect END_PROTECTED
