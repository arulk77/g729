`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFBTp7YK+wJ/FRkPBjGHSxkO/hdps3vUvsizX0Rs3lS0
ngn9w/TxNLwklch3VTYNnhjcD1fLz4Y7AdSsersAhmHX9x5THJSohT1pDnb7F8A4
5QY9w6TvDIHAw0218LTG0v9yxHvNrsnfaa2FhQ7Ru2WUfof8IWoHERMi2MbzVXmv
WaeOwO/vRL2bfIAbEKXxIQL3X02s+oY+Z12+2b5EJERx+a1y8IlH2jMRoUv8Ng+k
JyLvrHEC0wtGKnxJOhctgIlrlUqKwuQKSsy14UmBZ8AYmIRirOa8z0lY9DSTnlIx
ZhsyDoN1IvcrCby/Sq7RBr+EI1WRqXXz1J66aTPnkHsMgMRjqFt04/q/wMbs/Udk
9ILkWnMXzcCd0QtjK9yvf2Ut4TRpSa8pJnlWX/sdJ8tMa+Wmpv0JoToqoEoD0exw
cSJLPiKnH/jb9/z6Zef+Og==
`protect END_PROTECTED
