`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41gi+bNFADRD7GHT8eCTlmbXNPaJYHwbE1DDm6LhUSZZ
SlkN8HaL+rojGoYnD68eTQ7SijezTyhyJBts+6J93qbaQDzLZtJRCBAct55Wg2Ll
vF5QvtVNLHYpuNegTnbYviKBQWzEEaSD0nTrgKHifPvM8xsNb/GMbHoFM3xYgQLQ
sUoXv24TesqPQ5xpweiRbIO/qCAIcSoM7O0iYju9efZZraZX+Ss6jJI1Os3rumyq
SuXoT78BvnkXZHpqDkxPmppazJ40cxlkNBW9j80f0LyTrq08nhDg59wtrBmkk1XK
dm9A4cH4tmGvzDnAeP9rmg==
`protect END_PROTECTED
