`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48bzHbydhV9wDTvOtN7esxQv34/7wxHnNFMe02HTQf0R
L+Kn0AEGdHsx4o47QOlXKq3acrDm6+4Ve/pK836h68TOeiy1SMi9eh9GrGwAw/AV
Qd3n1Kp6uTL7BJ238lz57t33pzu3UTfijmxRXpRuJ77BXYLw8PPdQ4iX2webhDqc
FGsE/kz9P/mdasjSjgwikQ==
`protect END_PROTECTED
