`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBsNl9uvvueg/1DTxLFBXhTzeXQSrL0C/M4Gn8KgZqJe
5EObXBCU+U72/7fZD+EVEptNlZwFOf0TfWZCt1Nu8ADmP1+j5yxqo3eRCSXKG5mD
TgEdoADMjunE6Dj4+w5X8N78GSLZEz/2TSzYaf7BDJt78Skw+4sNzCOKFTluwj3d
IFPeG5aOKB5X2iH1HLNs6veodwscwlTqXeyHLdRkS9iUe2McgIWQa73je/Ht6ZYf
vGsk+vRHR6/W9fzlk3Mm3ZOGyeaxl5FV1Yn/Yru7dX9fQiK2SmMLo+ARf2CB5pKg
C/T9LfChHIHvRofxxvNdm+oAhLFkCHrUABteftmYMu3HX6cJEcdlTUXetBvdyAbw
b1WJU4EVFM8nln5cHKc6Og==
`protect END_PROTECTED
