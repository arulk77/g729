`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCny6OHXG1ueRvhHcQNGqTs6hWonJ3q65YDZFHe1yXOD
u63IUAIfyjhb2F4kMVw6qjt1T2gNfIxZP2FuIo1fmlzGCc/armRdkHqlkX9N+rh7
ElDhxr6rOoSlYzqywfmnZrPOrU7TYkg651wr6+Q0p/wUp7jvDJfH6I+qtrZIgjCH
22c8nvGY23TUz3clSRb8QRPBC3HUPDCGnIsAovsV3U0erNPDZYFS+sbb/35OfAsE
yMwhIe1xObDLlWXwIgI6sNGCayxLQxe+fvTRz+cJPW04JbA/47NMejAOpL9ul8bS
xggFcrqSS/aUtb60u5TUNe5o0rKP7Z6uFmPlrtqx8VlhzUXOombiHfP2BOgQLi6x
LPXt6cbxq8umXY7lvrS1sikCirrm0HKlbzrb8E9CJz9y3fVB3DV5qODBcAO4Jufj
m2lx5y2QEGNud/Y33jgHZIxBwFVG7RjaH/WXyx+DJvpCaDqM4Ipl36eqMV7WIUjq
LhD+n6l2FY8K+KV8Sbp/OM+euDjTKkEsHGhiFWCB1rftt1jhuJY+55byFxNqkcCv
I24BV+xove1Q93sS7nGZJEJIIlxWuQNHfumz/xpurZMO2tITJSDtN4rQ3xU9aRBo
+EWcdSmplSN+aezuD9jULtpcH9d5WaguKYOKJLSrFCAqElHILXN//vA5gsIY8hB3
`protect END_PROTECTED
