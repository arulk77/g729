`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL/3HzXmriK3buWPCZQIF+GH7gBRYT93OKboUfhfsjJK
+mUQhstF+94W1ZGTfvoeLJ4ksF3cWranGpsjx4Y4A8VICubcLRME9k6N2x0aI+v1
vx/5d8UD6dKmOoniGNo89VnZXq6Q3cHuahrUlhtVw0PZ2e6JO3VnuOs08t6f60Jt
Q5OfvSikYtUX1MprF8EfC9Om7yCSR5UIr0/CxtAKGNRG1O/RCYx0DWewu+Zs9GkV
Cjdsyca5iH7sPbHj0OYTYrDyzJGzKXfNmuNkBTImaLaqPLtS3EWJTODk1WYxzDem
TUWLwfg7FndA68iIa3SRpfkbZkKIATeuQWx+wqFG1QxYVCm0BJVsHEGcCG3SeGMu
UydynSasqTu9K8Z8MctBlE6Gf//WjU2APBI4X6PWtQ0qm4/KPoly8Jo3UWY3pHDp
BlVpsjVkRJO0paBpEA6LBmc13pIZ3YXNQRejFUipfbdh7vpe1T/NOC8455U6mJCO
l2K5pwAmtkWX2v4Pbd/sl+PXLDtSb5s+8hDRfSZhY70z+bJ6GqrOKMRm5c9tlAUd
`protect END_PROTECTED
