`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/SoiiISWgw3qQRtArKqgPTazjp7EiMPZvVxfPy2VNC3TYDL43g9/9KkmhCnHi5D0
j6jIcfImbQTql1n9TZ4J8JuZ7XxavW7/LMBEWo9QZpg3MNa1gcxOYMohKm0zsTOw
/RknoJg5Lof501fObalR9V8QRStsNAnKT5TNAcZ89PH3WvjmhSyr3l6rDaTwwPzr
yPXahbT+z9YTArVfQDDSAObTz1RvxTZ2HQF+PkyFrjNdbP2HoZhoUOED9csvu/vk
QBqB+Dyz1JjptSP2FJxWw7Ee7yJmIUZHminkKzQ+hRIQJ1y6JiyK+ap+SkmDoOiC
MY4LssFvdHisDpyw2PO5m8QxiMBfU6MoLSakbs6B/GgdEonCDbo+CIqdZ1crANZS
x9Dx2wn1wrGjGzSUnIcg+YzWvOXYslVoEO93ttoy2cWOLfuY+lrUv/KD4a+84QQs
ZdxRehtIUIHV/eGZ4MafNUqe5Lv9DHlc0CjLH9N+mei3CHFrDppRg+YtDvo+ri/G
uN8OO0KI7xzuxrzjJmq2GP+PJ2OqPR5wlh7aWO+mHm7NBE1wQzhzEVaz+fM29+GE
rnlIuJfo/bNrufe62yCraCQ8VDLyga6f6CKDsulRXp0q6aPm+yVvzqg2D/ZeVtiR
`protect END_PROTECTED
