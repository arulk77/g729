`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN34oWokV3DisogARRTS9n46xRjGkBe+skKSKQajgD0a
NOSlHUMbAWlj+JKLMT1iBa9T1c5KrRosr2xH2jyiWff1fSxUjRf/TIDpM9rz5MoL
dFBTEpoMQnCnNRoosFs0VTEF1+TrXSKopKOG6nLJJwDp3QTgZOSUmB3KR4t26FlA
7fmuJgDA8sXpZIKmR51sUaYGqY6uE1+I87gOPor0lJMSiSTwSP8IykR7811Qo35z
DtVGzOhdQq/B3w4GOcgQEwHmmZcqreKEqIa4qeKyoAKLJMLgTVKavUj6il2HO7+i
AqE2c7f/sRshdSNl/EV3IMOssx6hYVK/X2+WVQiM7U7TxbVC3XTpJz7d1/BDDaC/
k26OOys51ThV9aeqpwkuadWEzm1aqIU9FbXNGdYm1mPMgztrP5iJps13GM37IVEp
8QzTwMwcF+Y4k05lhRpqr2xe0QIeKj7JuqGyKG/CY/GqwNxSPJ8TCqvP1s/9mGhW
SMHNr8kZ9shYSHitijLeMA8tX9fgyczEkIfpNaoK4REy7tbaZCAqCqH2l+TkaP+f
FFy5+z6gEAujjD2+V4Opqu8GA5CendVQD59ofUpHVJp5wFeVcwNkTtsmbfKgh3PP
IVGTRpMUGKhlVVHblBlkNnI9s0z3SZx3Y3aENFzb1QTP7LUg/uOGu3Pk7dzp9eyX
8derG0kiFPCR30vRpw4VL81vCU1/Ylv9mZeuzmSknSxD4J9i8yeAxvrmgCJT58pZ
t6qH0wvSCxSh8txzMyFy995NzD4sCQTrxZEoZm4ryCuYr98xMXTumcSicUYrrWbt
9Pj4xb/QPRHlSlcH27MPOEGmMVBo9bVW86+Atp35HwRy1w5cqFJaGbvY9dMadaDy
nu0U1YLZeCrrYJLI2mc48+FLumMMNnwssEKOxBo2F0vc3qLgGaYQMnwL/Sspryxq
s1Guz0p8uweWDMdzX5h6kYzq713neR3oq816kXfZ77pIOIFqEGD2xvvYZ/Rl2I3D
oLu8am+cFoJRHng927EwsiR9/rBbvRqQf/nM+oJ0lQA5/UVBIZYHBgw9JX599nd1
d8qfMxBOYUGEH7sjQchkIcE/gmbQkiJZYWUnYQcaUz90u9Cs+Rs1+sK3AIvP8IaD
Z8P+Gx7dR28FWijX5V1WpBH3hVJ4lE09agt0xZZK6wBB9SXUhsUHZ9tXu+17WHoD
CIyqbwctsvtT4NPcGjFL6zh9ylumaPu16e0sb4Q/KvXJWeMLGMadNhvjiChmLDnb
`protect END_PROTECTED
