`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveESKBJrhd9eMoB49wj99yS6av/+OFeFt9KcV733T0u8R
5qnCfKrZYcdK0tOGuh8XKXnFJjKSONiT4FbGpKyWO1VyQFdsPrUYekGz7Hb4EV+h
MsUrWGVphWuSEeCb4Ql+lAHw1ZgDyyY48rwf79tjCz+cRjVkj/cDV7mDqAlNySVw
Uw24kugMrYgBY91cLzPT9XwTNLu2ZyOuRZ5dismv9+uIB9TR7JfDPuWs5a/GTma2
Fe/XDo+ZDD4lddLCuy/2yN01cOEWNMhiqbTob7LLSwr8581YMkscEBhuL52sV0OA
IJA9WoGxL0IgaefvGRDDZAgdwjszPzFU87gNeEQ6qBb6c2+x/7Wa1SIOSl+DR2+1
YQpd0ibIotWhs+tRLPs1Uo8AN43R/vsXOMtu7xPxOmoVFBhIHy2m9cO4IquHj2sA
kz3vHrvrexM4+hkRiQDKBRuti4Cz/YVeIyHnUmdAD32UMOlSxuwOZhbzz2uA5qGd
GflX1UBuqtv2HLaQFU2GeqYvehame5en3LpDyMnYWxZGt7dr3ERzvJPPKvwc7wzV
87jU/n1yqjrDGkr0GyIJzg==
`protect END_PROTECTED
