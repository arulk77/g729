`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIYEjqDK17VpYzvDxtP8B61gcQKq2Qxs2LC22XGGuSQl
k/N/7suIZUVcqyb9P/hXvn/FUFmvB7MojZT+shxao4mPoLDg6MpgP3rTaVtLGCvh
SU8baurdToe/j1ldM/QssDNGxa6OtOaT4SJ9NY2PvpBS02ZPtpP2WB6m6QGO9eX4
Jrw/RAO/vnB6R+YkC1zstGlbYJ+pcBrLLHNf+rFZJCsLpjAVHSYaVWl57w64atAl
`protect END_PROTECTED
