`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKDNzr/zF1I2TWVDU6QzKJA2qLK+gHo6KyunTj0mYWJD
QoxYupEhgaDHcei7cg2sAHAscZ7Db92bYwBDogkGb010PDchPc2+gHd1Xs6/u03s
LnbXXVmMd0Xl6foiNJehupFreJ5VKMr0H2/JVEpgv3EseL1y0ceKx2Ph+5ulsBS1
QtarhzwhFkQvNdqrBUzS1BkD+i1KsI0M5sAlWsbKTRfEwk6AkwxDePhKkjMfVr+6
iDx8rNiLaeNauiNbpD1bLuW2/8MbOV6j13LCBOVYZkdmlbGLYo2CAuFVKYk7AXXB
SHws51ItDy2gMtSuQ4dNGdSMYehM860k6yvM9CoYgX6GKmRZ/v6sZkUm3U/7xS2v
hD4Xb7FKIWeTe2hLg/PxkM3tVxL51rF+iMTbDRq2tv6cpNyXSIjQnStY54ATXsHt
xueLtyqO3Cpm6me41Hy7RJJXoIza8iP2UqQdYwWQ8XS5QhDdyXRXmbWf+BLzgpG0
4V0DVvQPQ63dfR8+9msmX1CDOJglAC78t+GgUaQWGEpKTuB+pcX90LLe5DuHnAxh
`protect END_PROTECTED
