`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0AmsuN/sAwxh6kCJ26jIwpB97Ze2dG/z08aIFnlY5arI2VIWmZ90G31/gStcsLX1
xMdjsKAVJ+Y++A1xeWe4gb/SkUwoQVEnUa92F4F4B0IAZeVSuxIQFNBQ9eachwBo
RvsowLCRBj3ecxMy2Yc/M7eYCB/2OK27H9qyhnTzJ2zqrU/YVw0dvb+UlFADQk9M
wQagLRj9oJ2QPWGAW85h5INNlTsCDAXemqD3pluhSeeJzqsiYvEduh7ENXfbhnxE
L17460hTyAg0om4k7488wsQiNIGBJ5XWsjcDs5tfHL4iM4ovAnVTQ6d18rqHR+M/
p75fBEihrmGnJmzQuD4L2NzDMn1Lie3rpUyBPiomC4c=
`protect END_PROTECTED
