`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBCNEkU0crFnVi6s3N6Kk5FvYMJhLNVzhlfWW/PUFgpe
9VbAFYDFbxhdAp7HPg5/t73KZKHJ9RbV0IvvDCyqnrqpxHAsfwqutleSeIMR4b+/
00OZteI7D9Yt1Zb70v6IYna9TZUE+RxtisX6eEjnZ8fdPRL22oqFefURjCVMmZKH
RlwtIVc8LjhssO1Ib9I/2PlLXDbevGL4E8dZlZQGfjpBPDcV5XjoB1czQtWzpRfW
pZavAhDktvy5iljTMI5EcVAj1RJK3fYHwX0s0w1hsBvNaxI/UmAc3/qwYBVwzh7T
skr4HniPDPgpS8zx2zUp+/RjDXqrWPBeKms/8myyI7p+Q/Xb5LGF74ZQc4Np55bW
1VDx3uCryJ8IyZnmNfQ8KkT7NJdoBa6Cys44XC/VDdFQJ1SVnkZZZKJBdAe+MHgw
w+vqKK1AHF+RG2j5/zDcUApNVX/HFfBTTxHD5UqJ2eB8C8w4MYluYhDBKsyrHwAn
rziYQIJohxJHi2BmrNo6d4OLDBjFh4yDhHSBwBb32pRBG53d7Uw9lBP0UCsv/CAC
ysVtc7fW+KN4tsMy4Vpg8HvB1SXdZkJfUvUaJHQ3hFkqsXPqx+URoMwfGqfa2V1S
JPpget3vJsVcxUR1sjkPUObroYf4uQq6/svZdeSnjSEp8fUSHk9ir1U8jwClR3Gm
LHgyct0Aii1yY1WFdWDZLJ95N7S2NtfPcVSEuwKqMamv3gkAwM4k719cntmQqVzD
vE1YmbbUeBy40WeYVKYtnyMCfd7LCdhe4mQVj7r0you4D9reNfHhZQB8y0gSvwGy
30Ij3aeoqsM2iUcD7lqk7Vg2a+BtpXACRUaTbKro4nIwVGhJ/hWPh7bUv0K4CPK6
jYGEy6wtSwtLxkRnyQF4yaNTH6VswcZASY2uakSmk8GFbU5/GkVf/04AVGanIPiz
r0q6PNOdH7xQSyE85DSC8R8svyP9OYbb8TytLgMMi3TSGD18DCsCbmnwnFNkOHaH
`protect END_PROTECTED
