`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGxBIeNFGcsVFgZnD/Un/Kv5k7KXTJhjofXIw99RNn8P
ZP9we8NX8+igxNySXguy96wxNJWLb8wjVHETTzbtvdpyJ/UgOkkp36Gmxol92762
QC2kWIjjJ+jv+o0YqEIuz8txIMlq/T3rhAwjDRNfU4Q2LLWr3E6bDtnPHvNubh84
QvWoh6KWlDm63jLjRRL/Lu1FCmYj8G+YmsC8AXhN0IFT5Ui7YNnW5sT5GPfpvuC6
`protect END_PROTECTED
