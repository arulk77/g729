`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49A/uKFhH0lZEFxG4tEMb6Vbuby8yatDb6u4xbzokyKk
XMLQOfY5rx9opy2zIrPDg5wgftUETXQDujT/VcwtqDBgixqQUHuFS9w8DHSZ0TN7
fCCjKJVqZWM6Ql2A1Kvwxdsq1xHkp89SpfWHke1t/S4G4Di9bdgzyuzbxRjNh8gL
YMpRk0V3P579B3BdhH7FWC1GAYRS6gSZ0FBj6GR0iab6czeNy1mUQWDvKMa/bKOk
FF/4ssGnPj7Ht6cdmleDjrb1g86ADZ87L4wJy004fnk=
`protect END_PROTECTED
