`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGi9ZDoUH2g1wxIajk7bdgbQDCnxluMWsrdoNxXUEizr
1+/EFcDrxQTLEmnD/W8Hxr29xK7wKojZcnc0UT1MHxODga2znGXcuouDR/FUL2Su
6paa7tGICKqJXmknV+V8XuzZ99ZVP/Kr+QCdP4dIGQjNaRESpiGR7bAeN2SGhBGL
yhUvcU6xW/uNT8fisSO8caUTcA1ovXNJ2hk5o5kVL7Ar12+MIvFXyeq0PRhb64Na
sGqMN0YuhRC6XPbZA7Lq52prbNpUFowdnO6SaZhUYIMm2tLff5Q1/o2cGt3XQDp+
JZwgqgCQ2F1pwJoB8K0MK8n11gmsNxwywKekhYarqZOOV0DQDUSfqwqHrLgv6I62
T4nxiq90PmJ9tnhHwxYkF4ig87MynzR/JOTsJcuBAabuErxH06UnB2eoAoYP4gGf
kRweiFyV0I0YmoLKu0buZO7OuaQbaihCIZMPU+5a4g0jp0JAGGlwO3lp1YrOSwUc
kdl9TkUOl7ezYjyWYEW5YUZv4t8N3qehid3gVKMmjoqL4EquQqw9XFEUpiCX1Ppq
`protect END_PROTECTED
