`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fy/yqtQg3dwTPyluz8LP+kSo53XH3tmQMg8Qun8iVmf0E/QBBMqkzFFwb1wtRSbU
Qz7mGwwblZfoRKC01gWbC1UMuTKx4FEWSG0Od8XLWKpsnZBbv7Vd3XjNRoTeKuBJ
EqVrFk3MpTR/hV6LDDJxKhvr2IMtljw8E5dqDc6DcztQPmWfpbv+qsQ3Oj3mGFAi
lLowp/Cc9AUDTbAKNLHKk+ixdFEsBLModyvrbsmTX/8=
`protect END_PROTECTED
