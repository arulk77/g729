`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMr0Vy3lOakSjIutmAanfz4w901LD7zZ6/gU2GecJgcj
NZrLndptkk7Ym0yGIkXdL2vSINnXzm8H04ENwwFBN65Fw8u9GtKasPFzvfK0sesA
QV4N2lQWYQWUAX6PSNgs5aczKoo8t847wxsjX/f/lYykCYHV0unobtFbMnAcYywr
1rvsa3rKVHlGHeBHohLuel+d3c/SmVow27AohgDAMhYjUesoFhpqCPIfwxx48YtW
Ja73ogax90XOOpiN07N4kUjL0DxAyhbttTDC1tIkvx1RAqZW+3qAgMNpPxEdbdZL
CByPvK0xgexMV3BrsusDeI4C57TUyROk3Ee3OgPpNOxhRLC60i3hHNeE+n/tSYRT
APj7D4vPQSqLhoLK/FU47ifNWMhmrllrcNm8qM+1cO3ula6Z6ofIxsdA5jRZSk0m
fClqWjzhVtkiauBmPFMxTx/cOlmuotB+BgGLMMCGXJLVoeYp7/kY9oNMGB7ZiUiZ
am860C91fRsDdCuTN3cITQAo+9R6UppjlyNZ+95uvUTS+AccJ0IVcMZ4xuT3mAEo
noRLlvUVGN/+RJkowaimtrlsmsQY52Ck0S/M0k/f+r+QjJSJk3oRlw11o/rDwk9S
7hl3i9HeBPLJHALuAVnB7Ly/NWX0yj5WrLGGncpr646/UjHT3gXgGYlnk3wMHHWW
`protect END_PROTECTED
