`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43Xqskbsd5gRlc6fswYgt+IHMQrwbUzMnEJCaeMxjOt6
9qRG0SSVkolDQyr2L0b/yT/IGGvkPyGXvz0PwCPJtC6MgxTUUJKZLcPamrKl/gFJ
hI/c6+X1rb4kkOX8yD58zMZRfhwlj4yHHTvAX++JNCft1sbHhs1cMQ2eDxMvAOHZ
jYqX14VoCjBpyHQXjvOtZIOZFatbjcFQ1ZrtlPyGBtjFrIr2DcBiF9gRZgmwIRWx
+WGVBFit2YWK1FtA+5QQ48PK9/OBn3IsYFTRIdl4HRI2mSd6cBFeMzfa/rWFGcvm
2thAp4O7hFK72EZ7wc9ymw==
`protect END_PROTECTED
