`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/TaLQDXC1iHXVPCEoDeNtJgw2OXfMCpHCV6p+Y/IsmDq
XbYvM1ShxJrdWMjCT17yAI7GE5E1Km20ejoTnjb5tKIovn46xe/NXpQu0QEmrLLb
ttKQoGLLhbDsHE10q+sHgiq5RooNkIauAemzpL+T9OjHk43o1Z2QLG8fuU/3VvXC
8O8A2wWj5vWSrA229ne41OhNkaZYdIlZvdzquxsx7Q2ETHtS8UyCSb9OPyn/UQFz
WT7ADnyTakUN8DM1HE3rkOjWoYUNAEe5irWMbjuNVrHAwfWBtl/5YT7itlxkfYmW
fafTUswCEpgedUlXPy/1FQrkJTw3hu2dnYNcNGH8mokKPcn/vOufJuIyBjlpR1x6
+AGhZFW8NpKhZwwf09Wt6RsQY+yx15arn6w2wXpIsnHNNS56oxzwGbMNsJbXxtJo
DoDQRYc2ZnbUjcx3oF26mZ1aSN0DDIxY1pE7lORKEtY=
`protect END_PROTECTED
