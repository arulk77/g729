`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46vuw3MuTsaf6yGSJKJW8f0zw37sXl4m+Dzp869CjQYZ
yO+258wat3MH/gEQtOsRxFaKXwMw/83HE4aWcxMjXmv4VZylxRTkki6hdsAyLZ48
WM49alUSCuSqxnY+Z619DvY5En1niGKSyVNLBcNXxNHWQhEKeT1UeWE6uC77TvhR
DlcyJHdiQ/EwIYXny8N7la6bzFMMnpnjdmsM/3QXjlE=
`protect END_PROTECTED
