`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveELRuZhXCvzt023Bep0RsVPjVeSkn/D5arGDFpJm3tav
0/svrMHJrvKt0rthVPSQoYdFF1Hv1tnxSd/OYJodXSYsEWbWGMolViu5WCU+iGhr
VjYTsWfDnCBSQ988QKdNfxJSOOfoieMnMWYguYQgGojlzwRzyrDD/OYKsh/4bBI0
qgLGEeOu5dwpSUqHEQA+8MkEafSNvxsi0fhVd+xlQ0pKjaISaZU02SVMlcLFumks
MjXbxDBBTIktPgJqRwMNT0kzTYyMMBkCUefJZXEd+PmNIa4Tk81prCthqggm5p49
uPFKmsjRuz6qM/nS8yZhg4m2oG/o+3raHiC9UzllhqSciagH6eMqCkdd5nYsQiAh
oDuhcMIripDVtPRXzlvcm7Nd4mC2+4fN3evTwT9JII17H9QcFX2ophmjThmgxNkH
OkR24T3dMlmZm+0xWypTe+n4kSFeuPizstpRxFWajPGGDItiq+Yc9yvjYJy285nu
SAL0/2B9JtqM48MBYiijz3O0gtUKjNzxHilMq32qTOHlCiI+NHIrwJ9S6oJ84n5H
boNNXapvHMAEr3piNtxyN2QIhOlGgsbnp+Zjmya4GRzLovHA8wNLoDhmib5VXDfz
tbDyK/RVvixY5LkC0Miu3j+DMoeSQTDoDNkjFrBokbKMvy6uiBZ0Gxw0eZoE/tsH
lYPxruzWFTDf3aTPw0IV3lPRMcV5oRIjfUzQDTSpya1XOcPFZZ/epU38aDno1RDw
RltNpJQv6JM10+DTsNJSUWrkNy/UPZSoQt3mRWfMIg0yZ3LCFPkfCCGDDP2tdULn
fP4hxo5720GSA31Yp0Rs6wiBmghuqr3eEg6Fx1teBKo=
`protect END_PROTECTED
