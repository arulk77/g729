`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveANUhqCnqimnGMeyucJVUE9SMv5+/k2s84QEoUhkLPFe
hb+/EDc7O5pQe2Jzc6Isx9LbATZmXRHrmjxBKYMvPYTw/uUCRogUVomTsxlpcD4M
G+uz/wsGL3OV48xIBN3c3jIAVe7MyR7E1aaUM+QxCkDMNzXc6guIkO/zN/QPOVmN
zcpLlEL0fN7Lgnmt5ALXAg==
`protect END_PROTECTED
