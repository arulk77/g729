library verilog;
use verilog.vl_types.all;
entity DSP48E is
    generic(
        SIM_MODE        : string  := "SAFE";
        ACASCREG        : integer := 1;
        ALUMODEREG      : integer := 1;
        AREG            : integer := 1;
        AUTORESET_PATTERN_DETECT: string  := "FALSE";
        AUTORESET_PATTERN_DETECT_OPTINV: string  := "MATCH";
        A_INPUT         : string  := "DIRECT";
        BCASCREG        : integer := 1;
        BREG            : integer := 1;
        B_INPUT         : string  := "DIRECT";
        CARRYINREG      : integer := 1;
        CARRYINSELREG   : integer := 1;
        CREG            : integer := 1;
      --MASK            : integer type with unrepresentable value!
        MREG            : integer := 1;
        MULTCARRYINREG  : integer := 1;
        OPMODEREG       : integer := 1;
        PATTERN         : integer := 0;
        PREG            : integer := 1;
        SEL_MASK        : string  := "MASK";
        SEL_PATTERN     : string  := "PATTERN";
        SEL_ROUNDING_MASK: string  := "SEL_MASK";
        USE_MULT        : string  := "MULT_S";
        USE_PATTERN_DETECT: string  := "NO_PATDET";
        USE_SIMD        : string  := "ONE48"
    );
    port(
        ACOUT           : out    vl_logic_vector(29 downto 0);
        BCOUT           : out    vl_logic_vector(17 downto 0);
        CARRYCASCOUT    : out    vl_logic;
        CARRYOUT        : out    vl_logic_vector(3 downto 0);
        MULTSIGNOUT     : out    vl_logic;
        OVERFLOW        : out    vl_logic;
        P               : out    vl_logic_vector(47 downto 0);
        PATTERNBDETECT  : out    vl_logic;
        PATTERNDETECT   : out    vl_logic;
        PCOUT           : out    vl_logic_vector(47 downto 0);
        UNDERFLOW       : out    vl_logic;
        A               : in     vl_logic_vector(29 downto 0);
        ACIN            : in     vl_logic_vector(29 downto 0);
        ALUMODE         : in     vl_logic_vector(3 downto 0);
        B               : in     vl_logic_vector(17 downto 0);
        BCIN            : in     vl_logic_vector(17 downto 0);
        C               : in     vl_logic_vector(47 downto 0);
        CARRYCASCIN     : in     vl_logic;
        CARRYIN         : in     vl_logic;
        CARRYINSEL      : in     vl_logic_vector(2 downto 0);
        CEA1            : in     vl_logic;
        CEA2            : in     vl_logic;
        CEALUMODE       : in     vl_logic;
        CEB1            : in     vl_logic;
        CEB2            : in     vl_logic;
        CEC             : in     vl_logic;
        CECARRYIN       : in     vl_logic;
        CECTRL          : in     vl_logic;
        CEM             : in     vl_logic;
        CEMULTCARRYIN   : in     vl_logic;
        CEP             : in     vl_logic;
        CLK             : in     vl_logic;
        MULTSIGNIN      : in     vl_logic;
        OPMODE          : in     vl_logic_vector(6 downto 0);
        PCIN            : in     vl_logic_vector(47 downto 0);
        RSTA            : in     vl_logic;
        RSTALLCARRYIN   : in     vl_logic;
        RSTALUMODE      : in     vl_logic;
        RSTB            : in     vl_logic;
        RSTC            : in     vl_logic;
        RSTCTRL         : in     vl_logic;
        RSTM            : in     vl_logic;
        RSTP            : in     vl_logic
    );
end DSP48E;
