`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEWk+TLMs7nIljMuCHA48YPRLVOzpK58G/1hIGwWY7A2
xgOAnbPt4cQaUrDm0kUUiz2t9DjSoGVx3L+ptEHOyPXwEAs4m+DLIE0AuTKMlfGS
zEl+U1DZcsNRfq8V1Qr1ewJI1wol/ecNWUzfW8SrstRc9a6hcrtiWlRBq4bZM4I/
s3K0fnxYAr/1BzihifEgW+33gUbTgDOMio7PxYd5CiWZfG3P7flCWItnVIECxQdj
9yYgQi686YzcoenaFxlF6w==
`protect END_PROTECTED
