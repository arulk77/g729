`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBXetgrYzvdJBoCeTarEu45Ho3fD09RxJ9TYzqntx9Fq
DAdPKZo+EVUXPNrU1io+XN5gc3J/O+BXk2E7ZaozVWS8gsjlACx4OHcKvU9uHHhF
H6ePefOhyIh2J2IWk6zAEYTkn7oR8adimmdPLYfA2wUl+RNIrclP6bzrHQCPGv9e
dj1VzAXdDgr+SI1R6G70sFhpTJ7qzSMGC/aeW3s46krW+XWcK5GvJwRF3St3w48L
CW8kfuhDsWQUQAJVx+WAeqd38tKf+Nlk/6Ap437NMOUl+/k2+6A61rPWJn341EMY
315jfVrlX5cpobNBuNhqM+c/ewqxYmR7OTyieK6zsO4d+Vz+I4JOVnY6BsxRRWAQ
FiumCrq4Dm45BU4eN3dh2nXPbWwyYtAfDc4MhzrH9gQLCHvWfyUuBcf/S8z+qeMD
G5OpfgK3RIyBaPfPJscdIAoTVilrfqSB1OAPWzwWrdamxF1tcFccOGE3pGQKEAkd
C7qCshvU7ZhuP6QeAhRngFeVAUYVEy9oIopnlipX4S6y0HZfsoR0WTpF4vQOOc2W
CuQXcspGcXWnm8mYQmJsztDE1Pkg+bFb67GJYzO3AoW0VyFeMBs5pvxJf0RdQ8S0
O7POI0+0jtLLrt/Svt3ug1eV8IL+3RqHEBHt0+uM378wWm9laPd9Gm+hUW76fJBU
i2FkVEbXHraUiLuenqSl6TxlMsttSsv/K0RXDRRaScFBeBqiAl2Hfb055/t3qVn+
vli9vxgWaVFRevcaG4LbbO5lDCzEhyr00Hv+N61r/oUPhZJnzspQUQqqNxCbxJGs
acQY6FVBCtePzRU2vsJSHZPDoxUCUoRYLJ5MYrPnrJs=
`protect END_PROTECTED
