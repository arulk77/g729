`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cMlyZgcvnjFf/vRqdowr3OjmBT+aYuqX/MKzziDikBwS
7BLAplqefW46hl6rXbNB0dKlXmL3Kt1pm5IjYtQLpPtsTr7zUAy42wrjQ7VDtXGY
X07Xh4O9Pk13pP1E/ULBHNdc5ypRk0LNn/8aE54CU+JZi9lE2ePZ6GU5x3ddOTQA
`protect END_PROTECTED
