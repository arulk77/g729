`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBT/bmWgjnYfgkRy7tU1G5wGgFOaQLBvzHlpp4ZYf8Eo
ccJ0Qji1B3Wno4o4flU8GmxW/JuDl0oNkuHCwzXDf3EgJbNFPaj6QZ/xuO39CNcw
MEdDbx+OiW8UfLI9WhA/a07YAVwbo8uxWhKNQoEdphUPkuaoYP0Effr8lte7nOt3
txaxSM7UYqWsXnbHvjLYMtKakGYLiBvTWiO0kb1WosbQNqiUZJVynDji0pLKGiUQ
cL7UochC7bQlWxhs/L0XDteqiZ6jUhBJoQWbBCK0/YqHIWLgoFwuY2OodGt6cfBq
qiJtRQCy87o3vhJfDnQCETsr0cxYike4OTS0NhC5l3qul50EC8IOo7tfqQh8kQ+Z
D/FcTWd0Z2TFbqmYinzytdmfnGnGZsqkWz1PDeh4iM7EFOWqR2ZTDcTDHm7h2vBx
JmBPLbEuJewStHjh+0YUTI2Z/LOmhzk/3Uz0LIUUPPzi/S6E2LOp/C+DHYj+ywvv
g0w93SktmpJ9VWGi5y1LeQQz2GkyIILUvB50BV99TUSUvLUff6fob9qx7EfsHnJu
LUlyxlPm9IBX7elUWsTGp8hmG5twO8W7qtrmyH7LohjPS2d1gHtajfqM3v0qvoYH
48CgwWCtjY10Kej8HAJW7LeWGvySlv5UdjdHqfx7DJmfNa6Oc4abmwVdWlGkuN2M
`protect END_PROTECTED
