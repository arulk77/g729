`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4dtWr0Y4x4YLKmMgF1kuXE3ghjGQP6gA6phuuDB/ZwxAy
xpaMYiLyPc4y5ClGSdI5NbTux68hz04WqDzaW2Qld0UfnHo4VCy3SCl5/2LWKC1H
4+6Sq5dGWHCesSL43hp2m+OMQ4l+C+sghHt9d1qAOmTeLokNMxRsKhZJAXF7vssp
`protect END_PROTECTED
