`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAfXOcDzzT672xOMcmJF72n7+sY7sDt0V8oHJraGUpkM
MW9+UYbr6h3GH/FPc8JA1srkZXcpIj0UUKyC3EaUDe0dt5f2Zwn/75zoKtr000bb
DLyOXejrJAbDMLR1OwSOHzI3Ze2EBUInYvZZuX02D8QJNb6eD5dnMkuiA5APZ62x
qR3H4S4vHbmNPy9dQ2ycSkEk3+ggHd4m3ghg4Fzb2Q9ee79jmjCk5/17MRkPdTGw
`protect END_PROTECTED
