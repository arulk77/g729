`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOzvHDInSNaMMkiCSn49W2rI7xUlaK+jYz4RgyuYAsLa
7VdeqAbUQU/fiY2NiaOl5FZXd/PVojo3/QzREU30+tlJSUjPW1z7861Pjyho/tVa
lTXiZvn7FsnyTlv93v5DUe+tuXTqQGO+yC7UNHofvGeQZ/yT6ilbnJVyljDNh6wI
zVYm45xiucOMlNpvi9Hv0/Xy0ynYqYBUlL7QIaviCQOlnhx8LTLhzg5J+GvPQR9G
qrCBCZ5ea0d9hjH0HEJFa0ULLv+MTmvH9C/15AEzyWvamVxRU3xt+85waTs4+JRt
nzdifTWlUSYoccColpk4MDUNau/vkqU/mL6sZyxZW98hEfmdS+MOcAFS2YONAasu
JzC9W5wX0izc25mI21at4LIL8NxwmIveOo7Kl/AnUTWpA8q072EeRjf1WTUphNWx
OUL7up2+wWClsCg0dKG8SJr+TN0DctUtSfyYRg9PEhxTtQAMsTsauT2eGFaZV7TF
1fscCGE9oGR4tjgIwKBzAkGL/HENGiOZUZiZPJ07CV/db1N+Z1JvJcDrMWKTtQdx
dWz+cmvJOrfHuDf8JmybO6SKqJe953g17EmJsHdUnn2R1bY5KwBH+SYdVM51XlgI
muRQczQpGrQIKMAMkSwKQBP88bOUsq8ZE3kW4ygOVAhQ/iNaJSXzvOF2R/4lzCK+
`protect END_PROTECTED
