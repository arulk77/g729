`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNMjodUGFjB0tgoFYUGgzY1Hz8FB8H1tyx8o8c6kuAhT
7VLUFJWEx5/kiRYw9ucEfyL44s2QS3Aoo9ls/6znxw20MvN8an4c80AAjsC/X2SW
1GuSYXhDgwNeq0fwbXvmdOJz4NZt68GXFfKPyAaQxVFy8AJaUZeAlamycJLQud6w
Mu96mNX0VgLV0z0eNgZr8HEHYPFS007fUk9MmjBcSC+iOnUjzA13zuvy89Ol8JhV
xNzxenJHtzF8r3QaqYvU19iku1r036qzlcOL9KRYJUPAcO9IVxhKhfIahaGy3476
7r9ZTxVeWC0AjJTv9E3joNEd4pMlcGSe5BzXptGoeUoShKpt+5GuVMwf2G7WsI5+
twG0hb6Ver0A4Hbf0P2dXeN9gJvrOSQNurZxdl3W1EtOItpPbCIThx3wX/ZW6NWG
BGCE+AW2rcUrj+TReyuwAw==
`protect END_PROTECTED
