`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9NKY9fOScleO8OQpTYNsYF7bH56EOq7d1meUPteDM309
DscCzGFXtU5CGDYSj8bzXiif6kFQOYXETJojaNo1KWh5KreHvn1UYz9HSoqaPem8
sy7nYNPtBQ+21moa/irqBFKMlvNZg7wNSCskZGo6iyMHRkYnDn/AL4wv+Sr4BBou
dWHZF8FWFKgQKls1YFNa+ReDzvtGVSGxrpMkY1YBN3g+KG1lR4VqLb2eNXJnq5G6
`protect END_PROTECTED
