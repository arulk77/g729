`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1acgb5369SaGGmClIf/GvEpyMGThROntZ9uPmT7McK7kE
CWeGdHBVPmi2ZiFuwRZ/oi/jizm/ZDeJJuVn03GihIu2SFD9PwDpXHmJ46lImuKB
XPFRYpdKjvSqnC8VFgwPjK9W8ESP8w5IPZizdfnCeKyz/tHb3DWxoIxXabLXBKey
QRZoeijaS+0tU8MmRcdtKtkAXD5giXoNV3VjdkCV27QX7TDimHBbirTxss2llZc0
`protect END_PROTECTED
