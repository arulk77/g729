`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49fNL8tWcCX1XHwdWPF1F8Llb8mG8zWyK3SHqJKInktz
mlJQj0jaEB7pc7BEsCe9VVXeejI6RzrYxzuW/p7tLLYt9Ay3Symf9T2n6KFiCeGS
xFrLUXDLV587NS+WXV5/ubtuj+kaVqaKMRNi4e76gy1l2O5oilfbLHst86wUghT0
pcCPPq53NZZATVL61MOcmJY/Oo3ETbOBTyVqooR5qydC9gJIHZR4rBwzES/2aMGL
Uk3JV/sIpCdAUP4n7w7nTXJZhCe4PNwhH/lglWbAKlBzrXbBw+N9UoCVkvAeeGBR
vueh2UTCPwtK9p6RqP+O8Q==
`protect END_PROTECTED
