`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLTzGhQE1+hsG0b6yDtEo4DoH9cyE3EIwuwX9SDEbrz1
mggzfTEn8uxjtU995X9QkJA4+z8u1TVleucBBFHO1l5wY5ivMmAh2hGZ2tG81IM/
6LRkmnP4i8ZlCWtlhvRo4s63xHD4VzRfkNg3wJyt/euqm5A+o9ND8YGCvGF5VD9U
`protect END_PROTECTED
