`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIbBa9q5JGAk1OARfbJiLWWHz9of8tXwVygpl6U+9snu
bMM6jtG6EJODeDmxN2R5bU7Ibo7cetgYaGRqtJ+nrBa1Zox6287AMfSNt/aTEsGM
kL61ebdA4pwc+BvcmQLJw9zXA4PtLFo2bZ5KWSQF9aO0447NHWY62n+hsEFJIAMB
XLxuO3V5Lj7oki3B4vA1d0Uukru+Hr37slh9eJrh1WcAwmogNAFeiSU/3pg5OY4I
qdzAvZEJ0LXiwJ/0tPGlMsn7eF2nxiTkPJjnjNzcmoG+stVALq56uEEUJ3NL03ge
bvtYK22LRIlMvUFgiJg5R6xcUhmuyOkQeQGOr4t5f7T2Z6c+rvgwilyah0vEhEUh
060jwShK/uqWMhWtnLSVCSySh3IHi8AYwQnxrCr/a4yVamJashXdYA1lwVN0PQDM
30Xrqgop88EBnI78pt6qZgt/XgLZIdImSToHFGlufbQ=
`protect END_PROTECTED
