`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHny+AAVD15TKIgprBTcnclbWbIgdwvtRt/tTArTJmcK
8y/7jM8wVKt/O/l0/wNygAiqJOhotYttDvgbNGUum43PY+N/QCM/H+lYfk5xojJs
MG0GIoS+kY+PcUUGiq4ZQC7OuGSr0juPDlPO3IptuTzmS6178WLelf2ND+VE+QlN
swRCfCZpdafgwXkpP/xLAisMaaKukKOehdNXqPgpjE0c7/R54kMt9e/nlTrvz8VT
`protect END_PROTECTED
