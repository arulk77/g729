`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOyHfW5HkoEVS+mfdPxAo+PvX89wQ8WxLzElabHV9bIk
TMAUzIo+LoP3SE1PzvnSmKCaXWSuJ8AmFWjPFJSY9l/oTWBraihRFTzVgEjQF/wg
GBIkf9PbGorFjHT1ra9UPs1U2gALgE4nYRu4zvqTP8eabScidVpjZF59lvjLXo7B
FoV39D9J2hZv4QdFEGleWs9TKFbLJAw/2VVGWSsKdz6yEXc3FMbcbMTKNqVpCXkw
`protect END_PROTECTED
