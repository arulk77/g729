`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
07xova/q+c4w19xa5tzWnutmQDy879BO5tSBqVaPPJ70wIXsXHQBMnNKgmSH2qeL
lsiezanQ9eS+Gyn0b8CLhSue/WyOTV5RMW/ogK7UG74sJJVDK098Jpln75nmFTDC
nROGtVYisYDTU3ArSdmkrZmZd+iHiqannT+NErZFqFK1swbVYPrn1CSNu7EjM4W4
TnCUfvzrGSu9H/7wL3TzoEP51wG6DllZ/z5EiWVrew4=
`protect END_PROTECTED
