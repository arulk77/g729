`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLfYfEUnE/xIYBmRIFjxZqGGly8R/yQbD7u/c2mRZkva
Nwd29Oqr/renjWrLfqd82pjfflH4u/Nd5fDbloQzBOoGLjtfsXMYzgHOD623M8Uo
ApRXriqxIR+kKW8phPVAmqQv8+tonz4Guyg2Mk9eksIDixYt84TMc631qiIijLf0
1Fxxd+J6xRZT2Rh6k2bAq8aTDQlKA2erluAGCr1JEcELrCt1NqefdpePJNSvl7iy
`protect END_PROTECTED
