`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFtQ+0wIPKzUT9gJMTvb1QPSz/M6aAqg3/DKKwJ6Ca4N
RISS69BER3zpIWI3y+upPh+zewAyUK0HpOkXpsQQwE8+MaEmpolLR6o1u+MzlMzX
R2uftuvmIVqq074vjcLCFhJ5mQ0VubqZZGA4bgwNvz5l5H1mD2JRDNm0G3KhVx0Q
lpflxA4umAtI935eKn9MrEPhfVxlZue880lfsYnl9i2yB/H9uIG2gt/Cm8YPltso
gqH7uRbAjwF8UvxifoL2CjD1vmys/Rlz2HrghBaRcZEJrLUpxbesX201ZRM/zTk/
Rch0PzrMV0AugowjgX7EUKdTcBu+YMpte5JJvkhLUgjgTCzqDzUNj7l5AwDmJIep
knnSK3NIu1mQUazW1ShwCitvpKO9rRcGarI2k27HfpltAhqhaC0iD2gFf/JPF44J
7nXklXx74KgIvg5stWGS/JnCro5dLnqkdIzitnxUFWbMF5FK7Oi4BjEFuOkDD6mM
WgNUCtFl44ncZCV8iJ2v4Pu7gBEIym5t3P8XiUodb0NoS1+ODOBiojMCnt+IjRv5
DWfjUgo7xg7DTElmrNs+Y1VK0kkU3+zQepQZbn6QqMNq5T3ZSL8VD8ViQU8REh/7
`protect END_PROTECTED
