`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zWl2f99vszLfjjH7zueK3wKtiTy8cRq8153CEekaGWDLmTJHx+NH+x7owFkHEtr9
URVuxOZhOZ+UO6kVHNACehVLc2iRpIrCJ6Ssej4ItjJcUd7DjhqlKbchXd4H6AiU
pu97bzhI93FJw1b6kVHUs/xMAWyRMW5Gf8wRbm6M2l8kFnYZvCZ4auGMLG1RJ5jx
fQfU9SZhbM426X2+HKFTgHyGnLa+S91bvN5mwCAKh2y4XLKUaGWDq/4Nkg/Ef0nC
xhhj91KMkqTb6j4y/+3SS0hK2YeGn25QLfUfrMHNrTCT74DeXWWg+K/XaHgSWo10
4ahXuTPspAX5F3zeFb6UVigMAB7MttENMKdKjIFuTbk=
`protect END_PROTECTED
