`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PoHoZpQBuj3O71MEU3wFo4XkR8RrYoamTUIyz4DfvrBknOA2gNO3OZPCZHd8H5sy
JBxFOvCvum2enKw38uZEEKxjx0971taE4+AZc/GYjau/ps+iWcUOjQiyK+gt7cov
z5HVUbpmpjCJ2F8wdjAZAKT/OyAgOWH8vNcxYg4JX/hMvEusJHKVv+bOxk4ugWGP
StNjWmSUqTl4lzl9cLmNd50l2mkZC+32D4lp/ebUv97fO6ZdtZ7I9GVG8dfq0fch
VaeQQ1tUo3YRT3X5I+FTnyHmDJ2yyR6BGQewphO+8lRCoFNYNoHJwLqgIT3oFXLN
qE0rDn73FMmkxa+mMMvW/YL4UNa1ebYafc8NofddY6eyY/nIBn9c+ffIwkvJb5L/
mwRbCqxRquRvo6EBuy24wDz2u61OLJXiXW/+hVN6HYgWA0Zez+I/EM8bDnGThCAK
GihPymDtq/WaXn7Jfa6we/tfs5GJC9qGdEWD+z02VVbmXMa5vPeeVy5J10Dgb59G
bVz1aecIe8b+RVmyKiiaCJorb0Vlu/1tZZ10+7Vu2NwUv258Y0ZS2PgCbubfAGrs
tDX5qp7CBFtrR55fj5yGpBcLuHCj0yGm+96HJin6vVADDSf0cV+J6nW8vvioR2Mf
AfTwn1w+94RjbFNGx+ga+b9IHUv9n1eY1O/UU9gJvuETZEZBNQwF5mdn6Iof4oaK
Hof78paQT+srikgJu00qBNxdH4/dYTddCCDK5v6uFbLKk0MoW72YXVGiAJszJT52
TI/Pddg/hn/27x3I9Fmtf0G0WUboCzuUvVScx+i2s6eJTWs0sb0jPZE8rhOSO2xg
5LH/2lIoP9zo/o1ESdajXEMKP8iwALjDcwNTrRbu7ybPyIKt+iKD+U4vX1PTo+EE
IzW2uhdcwl7zwOlz/g3e0G3cB2b+DToBDooeNxSqSie13YPPwzzh8yvtKQOOHsNW
xM0MYJ0fXUJXYGX/mGoWhX37dJWkIN+T54yHPsYqy9EYbz150yexogkd1v3DgbCy
aU4t2EE699QVy2EHGv5o3jIqOyry1x5VE4PLxk0+qGKttWxN+GJVMPdCeA2Bsb/D
`protect END_PROTECTED
