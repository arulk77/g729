`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI8k9nCCUv2vfDtyg7tg5fvhENdOV1m6ThM3w5TGg2wb
RKy3nFbIjYKfefF19J3199ztfRtHycRvPLYRD36otpqlPofpMzvkY18R3pt/CyIJ
u8wL616NxxA3YzUvY31yqG+C5qf0rJehqP5eGfPQcgJ0esD+4iEivOPBlum7d8bs
34Gz/FpRNWz29WC+5vv9fzkxCedRV4Lb15U72doD/9aZc9EMW4Mifuj5KtYplTz7
SFWwEFEv+I0kbFr0Gkh1b+X7OZt5gfWAvsOcbngPzFCsXkXyM7Uvb2D0yUyQVMG7
KW1mv7+V/Vr2D7jbDT9srYayYtqZt4Ft/o9P8EvJkb+27heWjMGxgFnF6P7EDzyH
FV5NOPHIlmfxibw8ktjMPmG82+0yFmZhdxh8e1+MjhWRAOfnn8UepiIvAMnJJfiz
QFES49/UqCUD/xIPEtjAOO6zdxB2pDbnc4JE7tZnQYy8H6dB8iRFdnZi4emGW4im
`protect END_PROTECTED
