`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rXNfpPn2PYNqd9/j4lNAoWGX3uunYEPzP/a+lr7N0znGiKKZSziQhvWXm5+OVix4
NpxZzN4CASlDVjFn3Hj4C4b+UmKBE/4FNFYAd73C/V5X8EqEM1h6fLzQcmSfWRki
QpVsZKIn6nWg3AG6mUnXJtLklI27oIYPCUPa+Cci9w8Hd+PiIvHrX7yQ8p9/KACQ
gRj6pcZeGn6M4KuIpQFwBns7OrL9a1AX1zNn2ZF8I8Md3sWSAp8a90A0/ZnCxGEp
`protect END_PROTECTED
