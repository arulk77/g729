`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kJKFNfGgiADt4uwdMYFT9lf0vyDEWS7RO5uV1WqwElK5DR/KDudPIIXJvO1rtjEv
k2izcVeObidi20NjMCxv4T8/01yeNi9gpTKUeYL/Ud1+XOytNL3uYpVjVkH0RXCm
M2qQ+wVsMVgnZ9zsKFy7v85FDj64YJMB4b7CHVB3cZK3Pxi6ezb6O0swxSuQxOFc
1rqsV31ketbOgB+8x/BiC2HZvuTZrmyH2//MA8kzVgb9azhvlRL7HIVNAPFciKFR
H/p3c1pB6vtMx4d9FiTBwBRdw/Y2BkGjtxySW556tOd+evO4S4TAdLmlRi77iWmD
N1ChqE7C5rSDk/p456txPPVBTFFxVDOf7C4pJBYmX+s9LY3EOXOwc/ypnpnJiEOv
9yCZV5K1hDT0XiUOzsMU2hNNhukYmEWNbw7ZWiWD0s1Hz7nn6MzDo+9tWxHu6QS8
xD+ruuv3KaDmxii/H8Zob4UlzwT3fB/vQFga2StRzE79fDv/RRu3nz1XOjkcM4jK
bSO1Z0tHDRrw2sigeYPgIMuCx/EgL9q7aAf/UJ3zrOQX93maTRgJjFY66hnoyYrr
nagdpdyeI0DenEvq8XT7gjVjDNBaWeFzELi9uCSbiQU=
`protect END_PROTECTED
