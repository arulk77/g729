`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rkO3eAsbrQvbYbxDEtV0rTc9/LIrtojeR2QWm/1fZaCwYO24PTujYsLrpSN9v4+v
sQvHAbvIZAZXgEi4mNdYJujfh9Q/3pdZXV7Y0cXv11K5QlLgvw9enZd6uqMyceir
ztAcWKW/crAgbVccHXkys3ZPS2G652B1X9vH9liWs1G4asofAR4KWj0JteF1YWwR
BkvPzmjjFK7YrdERo5/gGphioevI0lWCPoJMbwB6FIo++ud+n6Q0TL0xFx5d1+EF
4oSBlY5/gZ22NIYpUezpk86aivFkdHqs957scFgsCTChftWYH6BVSIduadDlJDFB
kCjasIcZhqbUMS01KmLcm3ah7a3DTQOf5eLD5WKjz9c=
`protect END_PROTECTED
