`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFX/uGx74whTrW4NQ+FMPq0F8XgCvBsBQACDso0DS0ml
gN3dXLODrHNsh2B7A55pnzQ5NnlJU7MAVOh5HU4O2sxoQOA4DJgIICL0XE1BTZMx
7Bu55PaNLWYuQoDL7RBKz/pElE0lXyqB10lbvRPokn0Y/aTT+DUyY+SLByuZiDjH
`protect END_PROTECTED
