`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
J8tIBe8g7ON5I219zEeuwtHTdHsr7rL3319TRYPllBktfMclc+GejhwTm1+uwdXZ
oLS4pTtePGdz90zm0KGY0iMeuBJH0N7rUxperyyE/5NqARpea1gwrj10X0+N0oX2
nyQ26iOSkdPNZ/JbnwT8QcOFpBMMVwbprdgyCiW0KK0Tijq+1H8R/Rhq+P00CoKu
oQEfCMRHWQlkBbguANrf9dg2C8lGqOFNTOSrE/qemqwooY7He0j/l5Kg5tUEu9ZV
pGa5X1PA94hviJprBSG+pHcpXEIwwXzPpOLkSIywSfEPJaYQsE3HOqLz9PPb7GN0
`protect END_PROTECTED
