`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFHuhm2z5dz486PhoP4idX7DFd09x6Hhboeo3HiET26n
gkf1V5eZ7n3Sy7cyeXK9ApHldnpfj33oKqMkxHLS9zpeGYw7yxmYU2d0uERKwbn4
quZIGUrs0BonlXPW6K4dWJLHMooH2ONdidDdJSVL5RZcVvQaWu5Yt14IeBd5ugfs
hh6X9j7tOS6ACGLhwfJfx9SakPw1WsOP/B34Mu2xPmHJyQl3W+8DjiCt/BPG3URO
Wr1XLj1Hsf26ceQeodDrXw==
`protect END_PROTECTED
