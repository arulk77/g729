`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/y76CQyNFQMY2IwI/MlBUmAB3h0kKLM51NySTdK76XVQXD58pCXiDq3i33z6gCd9
iZRK+BtLxYl6e5Tbhjw0bJDxARlxYsuDmXo1HeK2LlsypbyisRFP84agq0ezP/Sg
YaaITrVAjetm6PZ6Olw64G8CDxfj12Qtr/RTq1UqDAXkPdFU+wqVGU6LhVTeJIVM
SSn33SJdcZa18pHiXivVgtQ0hrFKFslRZl3AYcuh7yRSY7ZHVvvRed54AEaE5FAE
NMe0q86UQlRHKQRUaklVNFnNN4Gx0rG0qVhwsrYQ1Pfu9RQlejznphmTKGIS2nCg
71q8/WDIyzLiEJK0Smb+FY8SZhCqSvw2jx084S7g/CvYtcnGF8K5EdwjjjDPky6I
FvkacuOhcVMMFQSFlWHE6d+r+C7DEuLLn0Gz5cqzKCsAx33il6F6iD9xMPHM/2pL
j3kQpdRHUlhUfcQ/Uos2sLL3D1C3sNuVB3qXAuq2LeM=
`protect END_PROTECTED
