`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1ac9b3r/f+lOrHPuFChyhZeZtx9Z0+b25fBtkDaOKssnt
IEyJc5RZ9iRIgGqUQGPO3harziFdwrjCI9+J0aNhd8a9fntS9PaOzAohVnswz9cf
77VtOE6lQufZ5R7MST+8w0fNa51JQP6kYaYJovZ+cuzO8nqOlvkB2/NHTepxwV4I
hRy73xKqso7FKcrPAvS7OtSJUqpT7ZJBU5OAJBhsz6whdQdIWDoeF6JZb7I7P/bz
`protect END_PROTECTED
