`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aae61GEe9BugMvsZ818z/mkAp1Nq46GkAsRxKhXLnqwQMcUWjVFbVLpa2rV3v9JZ
axCS3ySAvbFYLWqBwIopLZVWecoLHd8FiwFJObGbLbAyChZ/VJYfGmtH5WuDw6O7
S8TPjgr8HVS+qTdKo8CfGFdagjYZKIt9ahGiT+/0CIfv+F8WCtwYB69seWMZeKKM
YJHahSVUFPfVpZ0rs7zNnS8frts3ycY1iyxObvNMehWIHDUxNeXn/Vlz5E/17FBi
qyCn/rSuMYJ8KgITJ+v0107T3sGqGuIxVbGMrzXnr9XJKeHuDNJLMATlXP95VCdd
S3XSDNU5m7UvZexInyYPcsMRl3kWP3DCJfaZfTb2FkGLL0ffhmulQLX8lXHD4ci0
PKl584XBqKB/471zamA8+UhaAocpzgo6F3mNf4OSS+/N/P9L10OKGdGJR0iYs4su
vgzfcfWt/O95umbkLyV1/w85gDviq+53n/IcrwokX8XpRyvWljYykHsA57bWl77O
QksJCxK7g0J/RMPN3CsHZbG9Lj3PDgAkx5zRrKhZoSIeV6q1sZITD7cjoaZD7RV4
KxY4s699rLrlUrArHEo8pMY4P7osY8moYTKg/faqLR4p9WQs5zj+F3pd6+UjabRa
9pyRRmtlbbTX/wCFSRjeymhCrdezGIaoK91ZQhVahwbT6aqAfB2vGJcjNGhy37OK
4DIqmvRaf6vpZd4B69yFoyNqCMwkoGKrb5qsc6P35BmHV/dtqEmG+8sAk8bR0vIl
XfCPMeI9UX+6OlIFJ5fO9za78KaoNzzFWxYhhHcToOEoj8arriJnNxfv/R9Cyzfw
bMe8czsO8PA4Ml5oF+h4mg1+Tt6lfvQ+nT6M4PasyY1wcLuCgqA8+i4QgxgfvQ9x
kd2xUoNLuLr1Fb5O/F0xstLBBYR7JQmPxdgNRF9kMzlWMjMrHv7jTooJSjSAAzxu
fylrR1JehdqrIN93b3eP+VZaoJ2T0NtclN40Yc3x7gBwAmN5lfv8VHtzXEBwpah5
7ZgairDLfBM9GOMq+qUeBcA4MF1KJlQzobQQ13GW4j8dNrjfCe0uaDE8gdfs/18z
RFIbwm85kImSM7LeYE39g+EAURYRwgH10kH0PO8JrL21f4wCfsI4plYu1KNzyz82
7jvfQLG/HNBiTyjzeS6N8ZYXMrZYu8Hojw/6DUU3FG7jSlpfjn9bYnQG32Xr34Vo
0gRWxcFd/D+vKqDImLNbhr/EVtxOUdAYdcltI6l6LcyfQIkxyTW2Siwx9x8nN/pR
nNZQkSY3LqoKDbpngOxR4AhpQjAAXazSKBlyzGTCr0WVh2Z8c1dT8mWoxTmjZWz6
oDlDBR1615LPAc1Zl1sAwbzWBsWxYp48NnA9f73itVCq9NubIrCYiYyroFY07td3
ECyeEDqG3kAtRXs6saIb1Xc52SM72yj7v6XjffublmWwHIocnXLMHlrDFUHZnbKp
fxcwpjB+/x5auucAEdCTp/fwCq62NoK1F8vkchyfNNm2cXb5y58hMyeFsEy5dAyO
/4bHHRQzuOp5D0MoKqr+LDgwCMugvUSLcgt5aHVzJwCHhhWBfU6WJKJEL+QOUaja
KjojO5voReeNdskozCc+4NGFm440spKDISgu+GQW6Yk2KVh3OmAUoSt60C1c+YNC
QSQfHsZNo7Cm8m3OBm8P1A6+XIgccPbGhEvaWwSumrUIsSRvadamg87plbajhfjh
Jo98FTOLvVeXeh37CqEY0wLcOkct989LcNdWLpswqsMOeiKvIV3sbwBzhs8X+9e3
t/WgsoR053aB5gDHwgT//2XMrDKtP8JeACHkmZUzJbAUHMmd7X30Uryczzq5p5dh
f8EXEnlAMu8eWu1SXb7sVVsWLvfCHHm9WwE4CY16oMJwl20DD8/O8HK6Kd+KuLgM
0CWRjoliar3hgPefgR6+WA==
`protect END_PROTECTED
