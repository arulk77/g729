`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDRPe8JaYnvWykzGsfsoiDmmOr294hrOY+Lox0gWGN//
y3/+gZAjOpw+yQDWYburmJvJHKWJZsyOqL0XIX71QZ021Z4egpqF9EBC7lzxcm2W
vUMXcH/qFEaXaIc607relrqb9AbYqu0zQ7jDxNhfcCe4phvsckzs3lFUdSloSizI
WRPQUA5rsvGeZX5JbdIteG3MMC8t88vpjIFv/dxEUioOb+f3jZyUB2KFQ2Jl2GrB
lKlrqVhfQ3z4j3CPSIl1kU+kYlkaJnKBoVKBGvTByi47FBRXM9NBaNgFldwlTDyG
xoBo6drE4C8GJDDOeWY2LlS7UQoyRtFWxa/HfKN3d0c=
`protect END_PROTECTED
