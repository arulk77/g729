`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43nNYy7eEVbL+b2Ol9zH2Pg20T24+o+RMXrfuweJOir7
ZT4EkJVpKLINr6N6kV9EIsGaG0jzR214YQlaUL9hIe62KxgC4ORTMzBXZTZcxeDN
8cuZLEdwwAhR3jHX2qdEW+uapsGB89aF5D6WsBw2d83RazPDCjJYq/C8tbGa2hEu
3dc+UCWLFODZu70vQEouSfVxrqA+0CG+TFCly6WCfH4=
`protect END_PROTECTED
