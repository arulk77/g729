`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41hgCHG7e6eBonMWq9FMJoo70Cqe9cZQ8rYvzxoY91LH
k+UbhkUqlpyDLQTc08orM9WU8kAEgGAVRm8GLNrYJXn0mfV+egRI7LwmYTe9aEQj
f7QY2idUFCtItFkNv5sVLyFoaFLSmQoUlsPQy4RPsuKyvOXCkpaKBRuse0t7k8Dk
4sRvzLGiWR6aLIzS+yhM58emFadhZJNZlEHF6dWg94z1Sq9XAy8vt6qruLJAMYsT
U0EQhkuxRgqxqnr8lDLh90wOksNr7WS2MJo9XbIqwKA=
`protect END_PROTECTED
