`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48glia4tM7kdqTTgZUDk5m5CW6a0LASRHyprv24EgSHm
IUypduZMUNWFVbZ4RSOgPGWG1MTP0R5+njZrhX8S8Lr6Mq0zKkzfAzw2jVWpFl2Y
hQjWsrzF0dTBfZECptx6qJcBlHGRPLq4K9cJ2XY5r68gGWy56D4ixCopRPwg3Iss
YRuclgnAb4ppx7In7Xcw4tegpcwdETqp5kEx91dIhoNxou0FGr4UEcfHPY8o7ZCy
waZ+XNJ+9ay264kKYkAghOm0kDAdYMkodEpwS1ynzo49XfwMsdozFplV/DCTeDez
i7KG/2c0c+YSAUDAPUhtrh0XnofYmXQf+M5w9Ue9FwyPb5wF26avXNTBMQ/YIqPs
Id6bfm+tTL9pazAoTwjRRGUP8HNDG+/LIfvRIdaFZ8ftNhSo7QzXLEQATCWIGMql
nMveVNvSswwA5j24suEV3kGePTzbMfRj4oSbcSOkX/0oEfkS9DfIqEDqyCOPmWDN
afgyhcZDv5pVaBRyMC01AF52mPloog8u6szlU9tt5NVmJc4TenTCpO31aZh3mL9O
0QhXem4uQiFl8fajpijiKQmG1qPCGm5nV9y3gxJComZgfMdZD6s0khwqiNNhwQYQ
BU8LEiVLHpiWUjN+OYpdaDS3GkynjgzRrw4ZK4h9rCW3JDshdUggvjzrMmvsvYqC
TxtYHaQoLomDLW29sMy2UO4+a/VUNezojN2yxaROxrl/jOstw1oPTj55dh1NlAf0
+9av7lWH0Vb0gtax0yHrWkkjhAqL0B52jC6surhEmCbVZxHeBAi3groffMBZEWWm
JcIg001NJLiqHoj5tzXXEKOERkj5SJUsuvaI7T+OxDRPKEqq36fJxzNp4myW5jnI
asTG7xRNq+YLLG0uaMO1rA/ekZnPuxxcOHAvZ3v0OTCEtkXCyNlXqxFM2u9vlj6G
xfY83D2JClPxHSZfMhWe79yf+AdJ6o+Gz3boNOrq735h/UKnb2jVdLmmVv6WdEZR
S5HZ2HXv7u87gqMkSC1anSaljYoiHAIiX5YZ96yO1AyAN6plz/PyP/vYWRGBqRxO
N8SrlQu4G5bwNqbw+veCSNBTuXKJlMeQ/g/RMo2fb9JXaR4iPEOtizthJOBmjx6x
strNdCBcimZhcDCJfmvKr/SY0RuaZMhlhZojbYIiIRJf17ZahqHW7xoW6J625RgL
WIrXQjcrxaJuOrTEHd7yP6jx7pOZdDJMv8W1ndPmYuXNcheWEBU/GDQZXVtorWDU
imGGcBuH/Z+/SwVZxuGdJZ6NoR4mtnJd5bntEteljf6PXbblnukOegbLNUU3T1z/
m1FXQkR/VV2Zh2ip3Xw3Awrqey9reUIepY/i/BbVq1s9xOTAF9mG0GCXbSiuRtHD
SYU5LWTXzgz0t72nl7ErLzv7XGwThaQDqU3Ex1bjw7a7o/vxd7o4jjeJBbUtgO1J
17pGPFEa7omZ78nzg+4ujxKHGYZ8jXv3iNKRZSq82oxtyXwtiE9FM3D25jeuz5XM
RiWCwWmcZjzDTYFMYrHUzdNN0zAEX2esVSJxRQhhIJ44ksdO/DggrCX0PKTfMZN1
FBG7lIUOCOD/bmEHIRxQ7gEDZ6hf+2yx0xs+wvELhsplYbdE+wa2tMg+VNJzhQZt
dK7lLuV4NSwItRHCxekDQ6huH0wtpI4er0kF3fozP6aWFvu+Ng2gP0YXdxqS0WK/
AGyhNt/VDeS7QI0dpolb+jpDIDIOkyk9Bmt3PEyP53nFOgc2SgrsnQ8t6XlTgdYF
72U98ucuWLzaJp6QnpVnDzu5AOFHSMpgqKxIsB2Sesfi/ck/s84hrDp5yhMZNWsH
WTsSt9oXZ6hH9OnCzFJbpw4EuydRA6c70UiXOcmWjiFwE3Z6n7QOx+x94KVhxkLp
RF4Z1Uuuk+XxaYsH3j6fn7FlTh+JG4m1b8ZCdD3mWGv6gOducCBwhY9/R5MGyquw
HirmiV5dm9dgEELJwgsPX4uu9khY2Eo3rgoBlM7t8AyugvbvBJURj5XMspsDA7U6
B8dszQ6XQH72YTmlKZCAoLnIPTW9igIwjWYL3qKrkkGMXM+fC/OSFsI0N3pZVbPz
yqPnaSAg1Hdy9Yorx7O4cFsgbishVvDx4sMKmdk/wr/rnAXYQ/RKWTmBrvj6Ma7w
qTFORSD22AFWqykxBgFUzMX6UKatdXF9kSF2pIGz1ygQ1HMNdJvApCz545DZ18XK
T7pp9u9+6aB2xs8zp50U3/V7IqD6Ktly71+0c0TFRyWGzfU03DilLx5CV/x9W02S
5SaftZfN04mmcriJaSkF/51ksp+xwSfziwL6q4zKxTKXwqp6G6tBqhlQq7oT4n8a
+oIxw+x95fn0sSHV0JdTktcvBvjGTZW+10JF+F+Aduz+C9iTFQ0T466cZ4rnQ1cl
0YcPGktzjFYYKVfh+/uEc4n9o79/l2wrSkaosUfCtSWd1aW+oa+phlY5cxYXmhCk
tzUEa6PisdN52+wYoZZ8XezrZYKIQO9uf/uWNE8QgNfkZcMwOPcNfzh4UrQl4NY4
Ej2FBXDap3HLaNJKFK5xdu6trMzKuNqnKKelJx2N9MOKCAY7GZof/+j1R54EPeH4
t4U2H1YDl1O+kRSFcAPWI4JX12Y9dv/xyzIH1J79eMJQfDmyZK+cQXAjLuhwHseG
AhCJhD0OSFqA0ZHKR011EA4TMPoy6qnsAXPeKSJtgnF1ijGQVwYbi/m7UAc7CYfF
IPvB7E7OH1qh9F7tgppAXK07DLJxACdchczlcrTr+PU=
`protect END_PROTECTED
