`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41ateHvSkelNHE4qe0a8hWYi9lMr97HhXOdzyH/aDcCh
oWcBFKiNIAae0mSscOzMFAyeen68O1ys/CbcXmrBnaE6xkEan+uU6GNRLvgWQLJu
0DrcxGPijK8V4wHH/ODNFIEGXeNi6vIO4irpwIjCxu7J0Oai+rvRiSH4O/7OYPR1
O+9uZgLWmGCgsPijC+cOgQwx7a+MZtHZKcbdvTklyQw=
`protect END_PROTECTED
