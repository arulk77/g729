`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP5B0U6HZFITLeBvM3zbyo3hoZvplKL0UxvR5hiCHzP4
VzdePsx/bKX79DtsgkVFb5xKYE7fMjWoQ9zV5L+OT+vwcQ2ZwU7cHyHIt4yu/AuY
mu0GeQ/+gyXA6W1vEebDT5AXgV+0Rt7/DPZ4wfnpWRa8p/yaHYJ0iMkbUIG8vrA9
zSNzCbU4kEdH0AT4EEYCxw==
`protect END_PROTECTED
