`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40nAbbamvy9w1SR+bZ9cSJdYMHFaDwDh4jpUr+isr69U
smWKqhW/szBwgPr1z2Fp6ki0zIIKP5vbDcXN0fbwQ0OKZ+WsGGq95tvFk3FqXqTD
H3xqJtNASScXL/yqpTNbYJOh77diz4wCCPkUGHd9hnErrHu/qPWOaFfSVpPLe2xi
bdi9+zLKBJ56nZyQMRDT/q/DJSOe9IWC3vmVeHCZA0kHY2QZCqsPivH67CTlS5qp
cvT2Jt4v4uF49hLlypbWrBzH61dEFzMgvVPimTd4fKlbPs7alsIzAIYjCL0dvVzC
GgQzM4htYg0wA5/a3eEifnysypXI1mAzHH8FVgVEFfcdOJihURSfXvCrYBq71a6W
6NMwCR7OjDrEn3YxNEERiA==
`protect END_PROTECTED
