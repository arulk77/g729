`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDsah0ktzqPoAUhvbNz4dMfyePfdCGgL7TvWK4Uw4qZp
sC/O8lryYmEACR3SqqGBBr3V10IE44mBzH9ktb+D3VxtuiSdTnv9tLEHdq0sVah8
HLV6u/oVMf4fnZhgy+oLBme1F/85a9q62wsQnIgrhm1YZM4PHmfGqRgC39t9oVEK
qQzLrQS1tz+aPl1LkrnAQQCGxgIvwX5AeR3iAGvec29sdwGtlCcgZDQU8PHspSdz
1/blxUq1Oou8KXfCdbUqxg==
`protect END_PROTECTED
