`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD91Bfe91cXT78ZvobxG2gUiN5aIwL/Wn2sK8rwG2amf
ITI2ClLG1yloE7DAYw/KymvfuJWKxdCsJ9vGw5ZZHZiSV4pWTEk75Ay1JMdVqwXk
fhY6iNaGaXhGtfX4jce3/+41S7hODqheRjEpQGndvPBqZccXweIbG8r7iMRebzM0
SLamz0cHlikySL0TUWTI99wu2YMsnL1nd35iFPhR4+GhXBn+MRsF5lz2OR4KTssC
6VSuGRKf/oap8wzIanRVrfuWrF5kUt+L/uB8+3iHmPE1tKGzACqmiDV+ByAHFxag
ryr8leXABFZnzyt1ZafDsw==
`protect END_PROTECTED
