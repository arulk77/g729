`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOh+zO/1B2ImvtQWaoG/twmBoWKPYaYwe7XtJCbFWA0+
OZ3mtewcnwMPp49EKxkucw2u9k+egsxUEhlA90YIHsv2maa2VDpd7y8S3/l7YbJ7
l2R5+M17ewYWzqlwF9BRED4Ipk5KxicwtSJEWpA5WNQK5795fMtThqxuvS3z3XeA
2ZB/Ce0Seczi9MyDe22tZZ0/DngFqCW09zaasJbUHOwfMYS2PoIuIoj72DQEsNMX
KqxUlxir36xt7Gj1wcD4CCFQwPNI4SkvV1yG+YiwKhTHtyCzT13wyeD4gu6f5t3W
gwxiT2uUd1F3utQT2pX/aw==
`protect END_PROTECTED
