`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI2Tk+7gp6k9rJSymuGcU8Yx3Z3xQ6aEdfOGojzZQppm
2eayT1Nn5fUucFTy+sLjJB+kEcRxjSiISYs9x9oOwFiW9KJtEILP+qfkLQdlY/I2
JnIUgMLPmNgFGJ5uDO7uNtWBSuQjSnMqiHCgkDYf/6OxoJNpfzeAOwrE0RrY7sk9
v404RH51NT88O7l1QlPhDAV9r2ZhaeTxp4DlNXrKoFo1scpZSbAwWNKc+CiJ8UPr
`protect END_PROTECTED
