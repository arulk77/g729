`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJLmKaXOsAY51ein+vT1Vl0DV29fNM9mE+yhWSdZuHbl
qdWJQ6P0h39GJn8GLH+tzjJ5En+5EAsFjh2cKPK/b/qxCBVZ+fIBA4Lndiw7MU2z
S3ThA7LyFJye+cQxvRDqLm3FBqMNIxS2D30TK87aDgMqN00lrAmK4rlCfqr4lw3Z
Uc8t0//HNi2XEENzPO8QH0A/tcuhnZQ4Nzq0qniNT6JudcGppHOzcNldB57EnD/h
p9W8YLH48wAQlGoE83kEviQi/nFwr85yz06AMNySw6LgkftUOgSQyYVJPXq0/mXf
qSjC6bZFx2JvR/L5Rk5IUcXURvPKMI6JOzsUvctxUPTZ479ph/L6BlO3ZgEeiKZD
ngpF2lfi1Ik3YQZS41D+TEwXLFZpO4d3/n9sidDoILwS0gy3U4rBGIJVJ0yu9ZMu
Ds/lLZBUgsp31m/qhIRSCJPu4V6IL71GYHdqyYHMbNLOntros5Hhe2wlzUFfylTX
a+6ERkuiEcxjfB4hC3Fqgea4bWwsTybOIA91Y7bFkdr+gCoZ4Ta+LdE74o+LB6N8
yhPs2PdnzWO4tbH85NyuObyEUbU27b4bZMwX7x28P4kQz9VdSpc4+OM+8O1mxm3Y
`protect END_PROTECTED
