`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xVi71lTXNz0njcXZ0/NmPTQVFpmrMvcCOhcMKy9rRRO
hojkd04wu0ztxRspiVqokPMiHIIpl8pQ3QBIwyFy1HdKHUWvHYSiYliZ97ux0vMq
UshDWT40tQnYzVPjicL285I4OgWZiGhh2axt/6pWdKn+6221gg3TrGl3Cd9rLh34
2OExpixNt1TmnALL4EXOO88yKBRqukUana5qEMvSnbQLTjYrMawR50ezEZHGxVjF
UqAtxIXNQfZlk7ooli51ZVEr0eTVkp1hWkYBLqLNChbTwvdl5FEXFcJvMPN7y916
0OWo01qRecjMDiXFMU2Wtg==
`protect END_PROTECTED
