`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiK/vvdThR/4gvnGs6a62nS5WwNX3x7xW/7/pOEoGV7QAD
6b6ozOP+6fHZjipBiS68I0Cj9tveM81pXfvzhpz7XiuwmSLm2waJidrIjrjLCaSc
qFnsbL93biOj9zM9jOObL9K2cdogKUCxAopBdl6/mZ78rVQMp7jQOeV+JSnZCGMn
ayO45fl5mKrr1SAXazdRKQ==
`protect END_PROTECTED
