`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4y5LTdOOZTQbhWHpC1q4vLw8Cj9S2h0fz0MnqrPr+cod
KkXZmcKatU2gUR1zDfOQDn4JQ0E4gyybNDJ2zb99NPU8WzpIWjBjX42ztBYYwXNh
TGHsSkf69dgl2y6pVz6IeB89ON5qemZS7/bF+ERnjcK5NEg/WedQ4Sb/pq9yoH9K
M5Y6kp4FYhy5BBiome3cIiRk/qqea41BDWP1Ehu+Mu63IKb8XnOljyK/mZx+c8Hr
NeKUyRJK24tSItjglv/UqLE7BnXgXGBvi2zEAfpVXvLNoTW0M9EJCnuzeDjE9rsI
MjhepECpvPKbcLq/8KBZMFkKB/dAYlhoZJf8xhoVcUvJtM0OgPVZ07aNsRO9Hkd1
Vw1XLvOqR14gj7YPZhBUog==
`protect END_PROTECTED
