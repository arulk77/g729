`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bOEDozYVfDIzWyRUUoQzMDPJ1u22aQzZEpt8aQ1MWVm7rmZ4KcFFOOjAs4Cminky
xG3ywfQrSrY2qPzKExLFWe42Yt9EDG5QohwHrPBvEJn38MH99SfQ3uLKZeRc+qs/
xbW7Hi3s/0SVD+4dWPj/TfGKlA0ZvT6Ez1F4dfJuKqUHWU1eBGcjetHu5Xp5L/fD
`protect END_PROTECTED
