library verilog;
use verilog.vl_types.all;
entity RAMB8BWER is
    generic(
        DATA_WIDTH_A    : integer := 0;
        DATA_WIDTH_B    : integer := 0;
        DOA_REG         : integer := 0;
        DOB_REG         : integer := 0;
        EN_RSTRAM_A     : string  := "TRUE";
        EN_RSTRAM_B     : string  := "TRUE";
        INITP_00        : integer := 0;
        INITP_01        : integer := 0;
        INITP_02        : integer := 0;
        INITP_03        : integer := 0;
        INIT_00         : integer := 0;
        INIT_01         : integer := 0;
        INIT_02         : integer := 0;
        INIT_03         : integer := 0;
        INIT_04         : integer := 0;
        INIT_05         : integer := 0;
        INIT_06         : integer := 0;
        INIT_07         : integer := 0;
        INIT_08         : integer := 0;
        INIT_09         : integer := 0;
        INIT_0A         : integer := 0;
        INIT_0B         : integer := 0;
        INIT_0C         : integer := 0;
        INIT_0D         : integer := 0;
        INIT_0E         : integer := 0;
        INIT_0F         : integer := 0;
        INIT_10         : integer := 0;
        INIT_11         : integer := 0;
        INIT_12         : integer := 0;
        INIT_13         : integer := 0;
        INIT_14         : integer := 0;
        INIT_15         : integer := 0;
        INIT_16         : integer := 0;
        INIT_17         : integer := 0;
        INIT_18         : integer := 0;
        INIT_19         : integer := 0;
        INIT_1A         : integer := 0;
        INIT_1B         : integer := 0;
        INIT_1C         : integer := 0;
        INIT_1D         : integer := 0;
        INIT_1E         : integer := 0;
        INIT_1F         : integer := 0;
        INIT_A          : integer := 0;
        INIT_B          : integer := 0;
        INIT_FILE       : string  := "NONE";
        RAM_MODE        : string  := "TDP";
        RSTTYPE         : string  := "SYNC";
        RST_PRIORITY_A  : string  := "CE";
        RST_PRIORITY_B  : string  := "CE";
        SETUP_ALL       : integer := 1000;
        SETUP_READ_FIRST: integer := 3000;
        SIM_COLLISION_CHECK: string  := "ALL";
        SRVAL_A         : integer := 0;
        SRVAL_B         : integer := 0;
        WRITE_MODE_A    : string  := "WRITE_FIRST";
        WRITE_MODE_B    : string  := "WRITE_FIRST"
    );
    port(
        DOADO           : out    vl_logic_vector(15 downto 0);
        DOBDO           : out    vl_logic_vector(15 downto 0);
        DOPADOP         : out    vl_logic_vector(1 downto 0);
        DOPBDOP         : out    vl_logic_vector(1 downto 0);
        ADDRAWRADDR     : in     vl_logic_vector(12 downto 0);
        ADDRBRDADDR     : in     vl_logic_vector(12 downto 0);
        CLKAWRCLK       : in     vl_logic;
        CLKBRDCLK       : in     vl_logic;
        DIADI           : in     vl_logic_vector(15 downto 0);
        DIBDI           : in     vl_logic_vector(15 downto 0);
        DIPADIP         : in     vl_logic_vector(1 downto 0);
        DIPBDIP         : in     vl_logic_vector(1 downto 0);
        ENAWREN         : in     vl_logic;
        ENBRDEN         : in     vl_logic;
        REGCEA          : in     vl_logic;
        REGCEBREGCE     : in     vl_logic;
        RSTA            : in     vl_logic;
        RSTBRST         : in     vl_logic;
        WEAWEL          : in     vl_logic_vector(1 downto 0);
        WEBWEU          : in     vl_logic_vector(1 downto 0)
    );
end RAMB8BWER;
