`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+RwSEGomCYq2rfKZJ7gYtNC7b4PCbEa/9sjfEUWksMwWDTkOcF15LmImryfPlhgn
buYmbU4BNBu659ZCYrjZb1kkiFhN1cPKgjp2YDS0/swqWpcBvvrR6HO+n5GIK78R
y/aBZ/IIbkA+oNqyMNPrgyygP1Km/VCzydenlMCCxAL+tW6Qwu1Qv2YGy16BDEhW
n4H+8cYlEJ1hcU5W4BVr9M9pF9qHnFRP4ayfK0D5UJnvSLAdtHTjpYrnPxIeeVRt
xUk0pLDqDWiMl0D0nslC6nwp6jdUYlpl+vCMo5+Efxc=
`protect END_PROTECTED
