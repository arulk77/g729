`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQ0SNiMcJrl6gSbCyMzY1irbSkDjXS5aD8OxXPzKobqS
9OBKgyuK3pyx/0PDNxHSDyvyLdCSSSJ14+X6B1sAxkMO8KZLY+Lt6pCha1785C8X
0tZquebcN6YTVAMM2QB5xZs/oxv+tHO+2slefw4QHXscvaAMUJBdV/9CtFy8/R5H
BJkNCjlKzu8HbpJjFMiDvIDNy2ZkAI/IFmmC+ArBobohwljWeR3yQb2b6PYPnobX
O4UDjaeFZQv3NKdDOOibCSFmPx1nrKpP7y8LhEP093Hi8spFLy1C24u8OIyar1QR
6Wr7FtjUu5i7vixJicVfamsaEis3wuqNoanTBTNsg5nPwuFPIdA+bXWhCylaAkuJ
brnk+XKY3P6baliMwkLNje2L5rWTVRuCGRqHLgIXB1bSKs1LU4ueiWj10xB2G7pW
zgSiHXKA70v4wUyPh21JjTkdrIF0d908s4GqoBqbwoR64brpVj+YGhcBp074OOE5
E3f+JBlkJPZTAH8Mto7IKv/bDSZUT+D/w0uoE8cMPwtn8sAJ2l1T0OQ5fmGwhhTU
UjkaoEXoY0Eewzkac/YHi8vWdyj2NnOq/duSfmV/RkQdA9kHi9Lf/I5m+udBH+Ai
iPGjLxpN+p72j71cxS7vrxV/qO/mZ+LqDWG0hEmRJfDFLfOqZVdzFCogxaDbG3aS
axW6yBZi8/Ug6yxQoijazCPKuM5OC6eC6tm3bcbJiozMxgPup/h55nP6tS4kFRmk
VWq+df1SxJX/KZdwiZZ1AhJLTp/DrTkYhmwNvtorAykq805phqNybE8mGRzdNWa/
JfUQW5bfmU2sducNCnS10eyOfrya5mxCncWGKMtpAu8e9Unw74nDcXBF/QwlPojS
1Go0zydkr5Gt/cMvpAlnQv0lprrO6HkpXjWj/qUCiRBHCu1xghjXP9NWLLWTCyzD
SZhUhSyilsPW9oeCsa2NZnOj8/mI4ys7OjQY4JLvQRluLM9h228L52ngHxULUMLj
aWzaFbgMNeYRkdlyhJVlZhW8+Yk9ZtJ4SrNEcjQmvu3Cs130gYdo3jrvmgMmrTPY
SSniFIESrOs41LjeJ6K0TE59f49ViMI+SVx8tik8KMvmwMjw5sw0I7+ESvDXBmnA
KxSIc/IAS+h8BtaxHF4XXCoB4RBuxDZnhk90ONYocSZgF1ld06QUhoK7EtUD5KF3
exF9qd/M5hhksqLQZUXHXqZTE53ga5IxOkbjyURY6B/Xj6pYcjyrpxQKHsOx+cUF
6zOc0kkhLDbB1y1qccZvRziFQ+hyqs4HYGwgOnW0m2EBn0bvu9mq9YEL4C4YKdfY
UT1if4n8KHqGJ8inZgAy3uTNF/75sMOoUX2zMfL1YCaRDiu3nHYIjG+svpMLiQLC
Oq4gXCVr29Sihm2V578X7xcBRYUEDzLzN2/nCsF0R0oWbNPPRuGcJp7aoxzerL89
wY6RpleBs1+hTAs2KsUMPXE95+1L5wwAkYW7ospctmZkykU3LC+sopgay1s2oB8o
xN54j5NlXAq3JShT7d6nJHKUORyEF8Cag9zTvA/1aXoL9clzH/FnHiTCIACacHoZ
qF5zeOnDqCInGKHO0P0u9x6LeJdtlgYCz/uQszFGJBl6GyeQRjW2VGJuxByiAkZL
94pwMyDtpU5Bx4Vnh0CsymnZQQO15awL2TT0zAENCRGydX8XyHj96sY+Ab42DUCW
l9+chRj5lL0clJfyJhC5bHku3gPylZD8YZde7kK1EASgXaRBZGyryRpsgzbVp8Db
pi9MRcXdr7IsikqKkqe2D/dWA1vvot7S5f6JWzVIWNTzS5fd6+e77VQsxtCP3Hk5
3EX9kErYP7Fmo8Toj4y30NV8qR+Kimz8eSWEFrDSQvQOLc0WhQ+jjMtjGfw3wfoq
olhUeROPGxZbqCg/+cG1Hy3kZ0i8wEyW4NZj0GSgiJnVfEsoTCUa4k2syZTv+X2J
NC99lEldrd4Oj2Rn0ZkiR2LuDMtmPsFLgHNBYMjYcc6S74CQqXn54WsOopewcy8x
MYVOUZ/1qpKH2gZDiMj2SnszCTLT2+2iESvygBAy4MVn8g0smLdwhQsaYxJuZt2G
V2jd9JzjPFh3VUbLPa/M3o1oFX5smxTueJ11ZkGmOsSSfM5TJSygPiZed4snQJGy
+SVTNO700lfu/h46PVxvibKXycS06ZkQEGYLdnxkgxJo0mP3ypSx4T3mahzjQ0H/
Gmnc39Tz75yIPSp2ykboDd49FORjScE7VZXWDUIeHr2WPnhcS3INNuVOZeI/YO+k
Uj2lLrV9VZKWy83uoNI31CRJ9TH9xB7aWk6VKL+9YTc8ImEYE0Qc6C2GztoFQYeP
zJqCrkyP6Wyw/xzCcjnF7cR29FP9BPzLCb5QUkUtuABeLXGgDnPgvEx5qyfni7K4
K+Q5vWsPmJUtljlVb5HYK9Pts4I7L/UemjBTgc1udr4wZKF7dZ1wc1wKNQutGmqV
8tKCOHT9LUBK4w4WVu/VfLS6M85ldbVXhbj1G0k3r1dirGCWgWtzVGE8JCY5uEZN
7BJzv9KeQzr7GFdo8speQNWRmOUFr0ETHiuaUmxWvAZs8z7OcLpkSPVJW6RjeFCn
vSZaBaQ09eidK2N7aGcxdUzXZPVSqlx4REXLN7V5IQBk8cbDLOsPY9P3K+S1QV6S
ihfDVgwmN7mczaddBhD4//a8Seyi1RFUakZobpOcvRINuVqtGv7RdVhxGZe3QowI
EvBoMePNO/e9ZGiEt5Tz26hb1zGDsWyVwQ1t/iKVDvoHK2XVIRFewy0SsPK8NYgk
23MgKPAYyuN/y8fVoUoopleclhyD0d/HabTGD4LAGoYyuU2js4aEvVCH0GQwmnb2
md8ZZGvZDhD6iNm2Ev+X3AwhL31HcdxeOWokDhGPy86DgowQjRGIxjGSOHs82cUT
WewVNF/BCv9OcCR61VkluXASNb3iFxWKepd2LYq7dAbQyEHIXstYxSf+DHE1/L2e
jtK98n4O4SjJHi42FclMnmp9bijyWXk2MIo6hPAhceGTl/Ss3v3silixvnYOswm9
AJFKSfi/i6zTdKG7niP3zbsDOzmkMRZLWSPppxiVVzflzL9LCR+wI2VS+TyueU8e
MGFD/VQ3jC+EE/WfSN80er0nb6Yxx3WbYA5fn2Lc1gDWP08axjZdUF7i+BkiZ3/T
05yERVPHqpysiM1C9EOZIi9jKJOXzJnoiaQcvlTGPwN6UJmJbJaG7+ezcnZgjO7C
9XIrnenf8+EBqgS0VNCLlWJ3AFmEkQPVqpUPueZWNmbsYWUqQEDz7ZI8SCNL2u33
5p8klNwn77SQCrti06kobxW8rnlCy0e+gixYeDaYCmw5NQYpAaBfEwkqb3ohz7+s
Sp8hKRWc6vG905CGSW1ijIsoognJILRtNwnAvJIW4sRYvqs6/Bcj0QHtqVbka+jB
SBPQFau0rTCDwYP3Z4dssGDC9IS/en+OFEFFsr5H55cXZZpD5IwTnf47emwDc5N+
37K/m0P3W7WhhjjRyRcGpFj3G2cdqxTZTKrQaHVPwuywLB5IDPlzQbHTjy59iFd+
SSmu1REY6CtCtLC4WlmXQ+GzmqMcmCkb7EZQfl+UWCq6lr0Z0wNARkUcgeniW58B
e6ey3IFWnC4DqZQCk6L86FbvkhsOGJ0huY+YTIk/EsbBilMTSmp3yHe3DAqiQ4BW
pRRUuBbYhcfwQeipfg1CDUIymOYI3QZtXJYxkdpXB5P8tX24kmmzYjVWtQpeQ07c
uBiofefk89Rv8Nck0xBtlMS3CEbeEkDJ4S6ACIqPjBd+M9TyWuKFpe1F6yMr74HR
P6FZVgws2T3ZVs/nJkbKPN7W1orOPD84xKbvTbgMcugU1PBXAQl9WCY2yIrtV+vp
iTPpIs5yhbiharuN+/6lCEHlXzHCbe7A6ggdJFqdLknRgPK4maMVfI+aomZ9d6jA
uIGakgD90fIPpqWRQX1ZXo8ZJtL40ZNh8t3N9+QOWKY=
`protect END_PROTECTED
