`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RqMZUh6yJ2FCQ4uO9pHRSsX4a5Fu2g6/ECnFjZRNKhTeeX/YTtdxei99T63V5az6
QD/6Yxoef/EZm3LNSfgiy1d1wI7yPWQ5tcUFjdOF61eSrhxtm86RAhTuUVT4GmmT
5VVSHiC3Q0ey9QZIismo4seuHpi594D93RGaR8bSUNDkN5iZGstUg83lGQc7dAJc
7/QPRzu7wOYa+5c2rj57bWuH4v4cYl6rxK+0f1K63G5UATPyETZ3Dhy7K4wYi6O5
o0UTyj35KmcIgBzpn0nykCEWNOfdmUxLnp+5rW8o/b0=
`protect END_PROTECTED
