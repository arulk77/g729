`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHJVjgIihmPodMSAZ8x76UMZHZpOmGEnlrfojd9Q+fed
rja3d5E/O1ZTORdD81hWk+Oy8hcgKg3S2NgF8QUq74Z7HH59d+tb9UzCQyyf+rBE
D2CurA5V6jthz6aUluOvXMWIKzcT8dX6q915O2lsXOyPF4aIwIlwfqWrByLcksZH
OpoxNWUqbOhYGWRmcw7lz+jpEZgtKsKdjwqOHLf3AP3Hf8hYEG0EegTEa+6Nekyf
4sFtZ8COcemhaBc1o6GfUQ==
`protect END_PROTECTED
