`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIzRhgCntWP+U+mqo+xswyitvZOSu5UQCr8OoJch/1Cw
8idPN0adTTRdlE7MUlVPmr3O6tHFGi+1TUmwvqg2OXOmmfmYE/YXyBA7iuj0DUC4
rcPlrzY0w2cCuGrIh7GdwmW5UlPMvzEPsmsdKmj4CUz053Yu9ib+Hy4QyLmMZWBS
5RnZcjApJf1m0yaWSI74Ft0v6Q8CHScifpaiTs5o271nTtgv70Qb90tpw3c9q1If
DObGfQ+WOtVU32yATV2S3hb9U5hT0UNDxIKZJUWUeN4DFzO3h2sI3VJCd69a3Gyc
cMj/EQY5DjUV9IrfCobOWHDjI+Q9OQ5xy/Hel8C90VCjaWg35pmweVOPoiz7J/95
XXoCaJbTcs+/VuPJXHEcyEBzQbxdYV8in8MaO5CHGqHcq0lPZ4epVfDPmAD2OkZr
BwLBpEF+2V1e9XXlxFYQaQ==
`protect END_PROTECTED
