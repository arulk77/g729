`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNzcooPbzgBhD7pv1vHfmz8RhiCtD8M+UkzbrprwZFqn
G9uhyr9xJkaOqdRqvcQmj8zDUWxVxCvkqPGmN73oouQruq4/NY1IzGRk2x8eAjfp
4CXVgi5VUizBX8Cn/G8UAvSD16KY0ooOtUhAhb3nVKP8Mnzoe9dfyhhfg2Wm8RIm
xxusYChqbFgv6e1CNd94xcw9qc/yQMExWn9M4R8UDMftt0Sd0iBJ3k+c8Na1yqD9
ulD9x/yvOSqEC9Oc0obXMUmzLYEiW3Xx95KzLhuLYZsD4yrfXRZZj1H7agd/Xc88
d8YzROcMid+n1QJKOLqxHUuELmV9S+Y8FXriroSywqErHW/+G/4ulGnCsh6vCv/M
PXM3IEHA5VZX+7Lgr9ZCS9tzJ3Yye/5jTiNoQlRJBALDUaShpolTDU8KoR4dSycC
/pNeoO6NsczjffIQ6G8YPg==
`protect END_PROTECTED
