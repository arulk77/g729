`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF/rCcd7EYvcQZhTX6elg0zqQNx8Qc3C5nzpbQnJ9G1n
hSjUL876xDyiqJZqp8akULw85TM5tUsadWqpqD/TzmXhzrN0frJbCD0C+wWiHwXA
vR4SFlOtN+969fHe/ES70N2QGQcpANvlPDt4s9KoL5Xq4C9HkratfmC9DD9r3GOb
EsOltm472tWuOr+kSiJBfA==
`protect END_PROTECTED
