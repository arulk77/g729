`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ERSLGEtdtSc7odNh+K7sHj67N3C/TXewnFAV3AfvjjzuwXKda187KFJvjw4im/X5
hAtcxgkpR8NxTY2z9n33HoiNMNyirWVfYy/S1xb+h9fJjnMyK0XDw1J2GymzauaE
FP0uPHQeLF+TE1zgTX16KMM9goR0R+3wcvuABRoVKQxE8qjQ3QyFeC8RcBzJDoxa
YGEvkrDJzZRqLSRAtkO9lJIMaSQETdMWVqjaZo0WurbQjTo6G8GLGfZvbJ5YmKhz
GzcYNv+byXMvIqZ/JTMDCvb3K7tIj+7eLBFJW12fJp7r3okdrEf1tWJQEW5Tvx/e
0SdHr+1jHIngzsv5aCkbkVD+bBdVxucayiSZM1Mtk1+RYB2iISdeM1n93fYiD4gF
gJHEyNmqGi0VW1PV/jNgS8vveLa4ELeAcbdioBn8IXhDiivMjw2ihhBpptTEGswf
Gfvs9nkcjbMzSJDQfyHdRJORi2kQxInPJX/Q7B2oI1ueu6sevTnlMC+ZnOxR/1xc
DKALJEFDYtpUwoLQBdbC0hdN64SoHZ/kGTnH0wn2OjzqcpMVLt/44sW33+BpbvC/
W4pnKRlxr5hgtGKwLpiPQkuZY/YnLOy1wprymkXz0E7UUjaqnAtGLleNeAEaSQ12
CIV9ADDdpEs76BQgB31veCq+RYxVskbpJt5jd6b26pi6mkXJ53lQ3zKqGDoarko7
vlNGF3KhE3hA26N0Jop+kyr1QRXUs6Sx39hSGF4MDLPsYWgpdG76c+emnZ5ww6c2
BZpzMLTVkXcqcsLysMwz2RQShdyj50CSBVl6vjAAxATBCoJeP1ghkvzpLt/+5pg1
M7EM2B14QZQUC4BL3QaGONQK3Oa9NJ1FAnh335Zy+dJPJh1TCkBL88PfDrTQaWEJ
xhm7/MQZBq1PSnl2rKuKNvipv7PC3xWDn05U4f67WC0I4buXJpPDv8Y0skBxfblN
`protect END_PROTECTED
