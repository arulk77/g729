`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBnc8dTgWLShdMfUN2QPb6MlzQPbjwORMDTgPWiGWWZb
wj/lHyuN15kXGP0YEDiCHMcRD/T/rCagUko1QRiaw9Zj+ZQEEbSiMwKmnqu2N+x/
ePTi3NXA/20pDWcvctndi+w/PSkcCvAWQHQbqn9S7qaCKvbLj0muARzpCO+wZ0yD
ww739ngK92h4ns/0uzlZiuucSHyfBCN6k5Vth1X0ZpjLV6K5hro/YKTVuxvQ29Rn
HFs26pZE8UZHCbm6pFB6/rygJ4pxKKAFu4yYF40xIEeu9yRN7OwHCKOJ39pA3xya
RD1BM/82gZmRkdifa6E9Fw==
`protect END_PROTECTED
