`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDfOk2fTqrCRWjXAfa0s50Riyjql9PLqBxwTkyF6iocS
IuVwdRzbxoy25Z3aKbG6G5uZDHmVkvhpCv0iaei1S3MTLidpFIXEOdespQmWRaYT
uA/BkrQmDkHrTdN70FEL0pXnhYgb43iPPDqLjdQV+qLvGwUZLDOca2/niSTJXjXr
NlSnUV4H/jTFQw9OTNccEEv2UkrvDyDDxkzCl7OLRouItjlcTiLWQQBBEpSq29zZ
EuoHgKV2hmCk9s89cu8Qiv7wh1kds1tVuIPylvkIxe7seOFPLrz8qXtP5xWDRKNf
HZ4NmM0+iZ+qsq+pB7x8cNap8BJJBML9M6jn9Hrr8MC5Ku5EBF+hJTzRXeZ/JeIn
n7hAzvb0B0JF9YUjvR9D6g==
`protect END_PROTECTED
