`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMJqI8Qt5jwku6VKW2hya/8JReTvmq/1IAihnteQgUQh
XRadk9l7882Lb6OPgwf2S4HgKyXRACUPYyG02pMuc3XQEyKOtMz045bNjQ53jSo+
ybdFbJv7+m6Xne/tYMiq9dI4vXFFekVSItxTU298iSAEDaY49lLvCgMno1n4HR9e
a1FK0rr1pZL0MsiynzHdlCm6M04wunJFA/gWAm9J0KWDDsxaQmFUisgdlh7gNzqS
4Zj40EfjuuPGK7BXySriCoXrt8AJqWjrMueYsgVNofHTDby8LfNii/0JceaLQoYP
g2md0lF5TFJ2IfPDDqgJdkBprHRsNmB4DQCDg/B5u3qu5sJcTuW+htw9A8SyUJHm
Th333zLJE6IX7zTl5Y6nnXdt4ufl+Cpf6d4CKHfhFCoc16k6/pO4dh7CPZDpsRAO
eskQr5CIK0H/mGeDpj5XhA7BMG8EqqfAEHYceSpGdLeVq+54PuAACTvjSWf5IzGc
YUMPzhMfcpv8fFp0FM5DpB+2XA+XxOXFVdNIAF0TTRY4AxKr8Ezwki7JDA51BC/m
SF1VV+/g3ful3UBo7AHIHREckHT/skB2bITczDRX10SvvpyQRRW7iOimRRwpljRG
YWP+TzM0WXjq+0mAAmG9mmrrFjWCOcFXq2ZSWxEc5mnzNPi4yfyCoET9BYW1i0rl
8jmWAd3Yj2dEQ0BjabkMLw8Zy7UoPVuF+uzhC+xbX05GH1ijHjiAJcpKTrXxAh0f
6rdraLpgAovnSRGksxRYOV3JPHKFYzyGVPU9qw/Q2kek0/tYNMs6jZM80Rgxj5F1
m+YFjdp5XZ2VGZLagPT32zQzEDnhj2xuHwUxAAce0Me8bcUUZuSohqRZRMT8XD0p
pXnaMOOHTEFHLUqYk+UVsVjyevJ4sB9SflcxqBhobIAG1yFoLUQtnBBfbOMC2nj2
63kkK/0TfoDcv+eh+48lXvkPBVt+9aId4Mq+wRdmn+steUozA8e0HAnbIsIoZr4V
iz171tLLZkZk20cw8XZVQhGqfDLLISlgUXxAK3c9XsE/K7/xEo4Lj7X0LlaETaxz
kVJqdwPCrIMXxpSbZ4N3d4RbXEAmunOvuAROxkTSZ7P4z+Knmuboyd1/J59liYMl
0GZ0l7EcDYbUJdi+GWNALI2uNGwZP5If7BJJvox14v5X2GSGyibCFsB7AMPVfhnv
OqZaWsYVISg8CQ9o8F3jOXWIYsn59f+oWmWDg/vK3Q+wdBM9TBBUxk/591qEcuKj
clcMdBjTx3pdJ24Uovdt6k+5w46PlWcPxF3MYef8LhiQybyezQB2FG/q7ZB/vnGe
t/VLwyEJ8mEcSkIBBBusFf1svGjDY8narCWfmjTS4/MYYk8J0buXvZIp7O6zo3UZ
KudMRVgP3zQ8Ob4Tw1gmMHLJB/WCHKwLxmpZdQCivvu+Hpzlu7V5HiH/VzPJfuSR
KulLKT3l54Mvwev8uRCORq0WOjId9CWdDT0KJ6nFoTr/bK/Ii/98jUWNuzkRtuUU
cVTQHSWZrXsfMEVNyqtrwEHnbhRojjmByiznSlDiF6MDY+P5UBzNHfMzL0rKzyb/
LLB3JJNV+TWyuVN7T4rFIcXMYTS9+Fz8h9j20/NLxNCeC6xT6ZKIvzOG9u5hxZfB
ecJD6bVqEUNMBiMeU+Iep6KTfXqmrb4M8jbDhj6b1mz92+iKwGninanWlngksAxl
W6DP4yPUxHBKFMGwcS0g+n/xgv5ppWw4iW4ADLvW+Wu1H5muooVwU21iv+gzrzyJ
hud9veMGL+f3O9mMocP0dv5cl03ToU1hy8C3Fv2Cusuk0/S5u6PSTh4u9OO51j/n
2WMVxKiv/bSOxCkO8p3jk8BAt5ICstX8GS+P/8ilPpm7/epAGXjZwFg6VkHNi1N0
FPlqdGj9jaAz+nGOLGD1R6akhglCMpAZs3tL6uVMTHCjDgFurAM3RNKIoGunQz/x
6sXlS5Wl4/VR4bu5rfM4B4ivDdfG+o5l15QTMOCFkB7L9QLZWzAi7FZNzb5BTsbJ
B02UumAwd1Oke8MwlJd7MmLAhbMSjUsGcgugU++jAx2jzi86bNs4K9tynzAwL43g
G8hZK3/8C7SsZ8gBnN9E4TovwwsD+Wkgch+in3L+SZDTR2Ewcm/dsZSvnhMqCNZY
zAZlDhkWLU6vAg+WSuaKnUhLLX4X71FMkmZCqFe9hFAv5poLM58GFCmFUKDfc2ZD
h+26w3aoelpALsPwfxarlCpRKtDoK1jCL9/yT8kq2m5VgzcVZDBf2HTQu5yPTDT9
i27/lCN2XibxJkHNO8Kw8jkSWsXo/tDHE+vs49KqEIRqPI1LH7IYVV0ruWYwQf37
eN2Xs7YiJd6zdxqX8up/a1nOmmtjAT/acL8BPUzm7iSSKTA/LrRetoCgie0XpeGZ
ENvhicqJNmzDzuPnMlvLvSl7TMdmUKja9ZpMhtjg3qb1+hRYcIVxMzpAxlERkGc8
hXGhyBhgNWzOFIafTUWoo+ePUbqjzYJ7Ak3KlT/grwr2eJLrOwEXtqI49UslYBIZ
HTEZwvFG0xmz29hZJbopfos66islOkKXykRbcZSC6yrUMf39upXAgDXKgWxFhdGU
tFi6l8IVWTU75v93RjkJCk4ldGOiUQzQm0TAmQY8T5bc/4x0dBKPD8YnRfelT+WL
KimG02HJkEyTlJszUPJXU0DQNe8DbLhyNZj/KNyYFlUOPIBJaG5XG01H9ZFQx1BB
6zonKn3nkHl+NwzkdTPdUxAEPnyGdjONC1FFXdubjJazUxJOXNEikgKRi84JaaOq
c2Lr9zE5AxnzoKQojrtdS82vROEXKlboJcGUzugABbVXT6b7XtuB8ahuRLLkad7p
loIYl3Bt489D970kzs8vfgrPG94FSvpSMonojPJ+tZr8Dos5TBrzLRiIfmHqe2ey
IBoBfpy960zzU+yr9lYKqvpbX8o69M4/zoylcMSaiL0BgiayG7IhsrHWaeWRsUd2
2tIFsxOpTjw0tgFkL2L97EX8G0vmSn611Fmizu9zvsz3zBo7Qemr0MGkNTeuoURc
gErvxEEUl/xf0vUdKYZLJTFpVj5NDTZwpSvnhdi03hugFO3NGBfRmkavOKCZSO1m
DegJyz4ed4oRt7o76KUwatLjqtPRsguTaLoDM8fMbgokAssertsPlVGvwAydZOgG
6pd0vWFedy0VjrEmT0yrxaJ6bfspkDBq3uqNGhdmGpdoeyXOZp9WTSchOR40JQcP
0wtzhpTK2A2ECqqyQhJX4rjql3j6LWEsmGB3K0Gt/nqJHJtLfc75EJzs1FYpA6kG
GmqJQ+UaCJS+OPOF3/5bgqKRxUQrYnsk5HzzE/bEav5UE1hwBPSW+dSGkCvpQcDG
evfWAfTmbkNi8oOrv8toh4B4YGP2Hx2Gezk7GON2XMpYWAXc7a1NmNZ00/WO1mvX
XAzZU0kVuYTiR+PF8csdYDy3q01ElCzGlNehP2UFKyEGKjx4zMExcic2t0jhJ3dB
P0SepGhIDS2hRH1nj81jv8CRU27dbcnFu0m7rJkAhVrugU75NNukT5rk2IJzJUio
DPlkx947emdGAsHBli/rh/Ey2j3uUHiqCXheqZQWrtjj5i+ppizi7kyk24XPzTbw
nuI9mSMi5Bfl2/q7ihiY2gceo70ZqhkmWlWswOJR7ytQc+VM5fdyVuj8qPUu6jyX
i9gNKEq/kGDbhba9tVFee1NASZTGO9P2PEB2notc7q206QRUn5vqI+/htB2wk6QY
k2kE64/igVoTawsHSXGj+sgPdCougjfkX9rjC2wv8ClbqkaTKNHjRbhIihIXaPpK
sNw6iwxJc3OnVT+z9WtrD/ijz7YqJzdNHnGhYtytlMYThv9jeNMrh1dTPf3vZPkm
n6A02cenaXYHnubPHBRmLe9pYqJG2JSPx5DP4uuFxG//RyFAScSJ2dBHq6m79Vkx
y0wDJa121B/lPEQYk4+CG+UmCI+Guf4/dB7lFpKEgxgXN/go232PvqNCLcuhRieR
V7B7oqfUFP7ZTKoPjMOTxMc5lF3ntb+AkqnWuolpLy7C0GBy+5+9XVYsj1KBkLsU
YDJcL4HvtQfuuT8r087zswbDsI1XkpGRcBhmpWeFQMGDKOFbx9ncDEy9x1mLb5u0
bZSUcwVacacpxhOn2Ocy9k6aqs9xEMc9R3dgJVM7P9p2575t8HOCqXFc+1HOLLPh
AuAqaQPG5X7KxczDtkxT0rHdQYgQ0/CIaJfxSTNIHkVkBngh620GBIyUwrT7PcM8
xLqgZ2nZWzYjKpfnWGEmjlrXHNmRIW967vZNWKAxsvFOXVj8dL4DE6CgebCvf5KH
JFrOY5SyVQOzBLqhFqeBcm+7m0rZYrsXQvgJH6o+ehQIgTwH+RwSn2DFtTJhg0WY
uJRM2U8s93X02MJ0qijyFzMzJ+skNXfM8Y22p6o7SOF/svIAwdAcixHlQHliHtvn
oUbK0CfcTxS2Miy2rNoPiXpA1+qKB+yxDMFdb8z0VB2PEd/1vBi4b2c0B9pVb/Mu
1mZ3JTmT0cyRvjpG6TEz+spoCKdTDcSClGUoDLG531s=
`protect END_PROTECTED
