`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBK3qFp40n041QDDn8M2ypFoU0XCrqGQos68rG6XhN3/
UKZMz7paH9qL3akslWROn8RQBYb/3KwlzMOuHyJDdZkk48naf4oFkm4cK+C/KgBZ
aKgzVAamnRIDhplHTLng9ciwBCRatixJMZv5R1g0hfA+xPqEWCZMz7eNPUd0TzTv
1gQR6+t0xyNrVOL8y48jH85NSE4GGz36BiQZgXMn4xDqUgVi8yPl6aO463BHA1VM
4FHd2cvNdk6SP8ycctZkPNE81SWa/jJFFnM0+lRU+xevvFn8ZSCARt+n9xcwi8Wv
eEl4dBtACgshZDuJlWlhagVAc0UR5OuhKF3x9TrprAh3FpBIrZL+lzz8adOLtHmL
uCuSiYVT1XL1VmzMNP2E9GQJAGCcrjiPmlqsp/ZCtsMyZ0UAhTgnuydoQq919LBg
OzgEvUlAY308+eM30J+I7XEtgqaw04V0gMXT5E24RkNgFINxOB+aVi8GM4LqIDdd
wIVREeifdtFGRRPiHDD3WeE970548jfvVd54jiBf/fpqLGit781KCz3elyhjfQyI
3pcRXfJ6kkab4uz1ZpdTPOylBpeS1X+UNPtA2s8ncfo0Juk/5RRmHNaq/+y0NXX5
cV9n2atQuaeVPL3medD7bxK3LY46Et0HxQ+4fPip3sACZJRNtvvxtMyKd9Azza3j
dCEU/ilDVpqR9P7TmN1srF9tpov3gYq61Y1fo+eMnfPDJH7fOfznaqU00PRxJgVk
1ehjG4N4G32JwjAMxLdGYD4GTNPXbOVsmjrPbCfSe9lOZzGcHMs92aHoQtkw4LEC
SsrXGekRZprpLR/9dQBsDqfC6uUp2URymG4mx4p6WUyKZt61E0lcZzmJjP6Xnoty
ajKpiUeDOP8HTMObvV/QTOHH501z/of0GFMLV+22xzhQStwNeZyqnvhEe4tMgE/r
S/NgQxnja5lRmwalV1BnutfmKIVWEsuKh58PMbOp0oLd05yKc4ZSnGwcU1w5Qnxe
hoKzoWw3SItFYN6oHkirvDZYP2fNv+D3e09lbYlZ3IpG/ZSI+1R1pPS5JXCRA3O9
e+/ca0ttfO48QZUganVvwSh/WKacZOKTuTvzFXOSj5sxAIOQR9D0fcTqtHyXyZ0D
bidDHFqn+vppj8vLVRL0zvXpM0v4gf8GWqI7V5E4/PpifIqAPQKx+SzWhsiLElZ/
4jjzCYwrxPhMIUg5W86ffMCWVvW+j2QzA9YZjdOHnE8ZoQqmzUiOdLYqo0kefXoo
PxyZ11I9o+2wi1RHPzrKqEELA28weHWBSLu/EoApjb0s94Zky4kqdB/hWpTnbOLm
cyb4Wh2uKU+iy17GVMeXr9FvxXAXmbIoL5dtuJk/MbKkZhE9QuPAEtlsqBoao6jY
0gcQOIJAS+eeINZXVmGaWgDl+guT4XVP2/GPq0hCXjg0sphiGsd3Oep2+nc2C1J1
8O/sqO4rR+Xw3772qWL7XOaPbkpoArJn9wA5t4qd4cZkMF5QV28W9wr5JyUnaLpF
yS7ccNlsh6Pun8cjxuDGgLRSjmY+1i6onQ+yy6czhWTKMuoYh+6mvtEUnu4Lqouc
bfLL7YG+4V1vwdaqofuJtGKArREBjY+RnuhWQGYIWBE7HmGl5qA6N+hX6kNjt6xv
devnnRLCsj3KmKIZDku/uAqPM1ESmJQlgB1vP7hZXO/hrcf1TVV0LWiUFUkpAHd0
6oH8G2IuIv602Fw1DABKvwjeSUUHzzASU3nRvd7up0anEiAJSivtjIJ3YC4TVT+g
XPR8P2Orfu2DH4mcj13/SeRgwxqh4Ju6CxozJPdr75gosTgsoMOGhQpQ4F7yAVYL
/dzvugw8i+cSSYW0dQI3lJxo6brJKksatiy7Na2tnz4FDrEjj8lY7OrOqOGvkX2D
U83Ba+K5Z9DUtAQ/TdTrslrteZbkxbGTBxDwGUQXyD2oEKDciKxJzPUmGjce/hWU
Ip1OyxsojlAEfZjjMj3CayAls51cpE12M2iQu/9g2CpYaukQXJbFCnsPVyCPuVKN
DMvE31A/ZJWO8sX6FPeac6CmoFZ9hZypiGVLnIlfoMQdXd0aKORrE6g0fhsxF/cm
P72rindtTUSoATKDGd19BZ1x4kCnW96FpS4BPcnm7a9Jqp3EUu3Ogzbc7wCW4AAM
L9SPasxHlla/Sww1fATyvK0pH/NEBSn/XcBkVVcsLVPWXwjFUgj57nqDN4OEW7FY
woWEm44EeCj00fLSdXpkgiCAveVhkLxTbja1PchJJTlT9SIZ9ROgVdLAVrFtlgzV
3kjiTt4jr/wu2DZfi+NSCoJE5192DMV6gjrtIfivCsu4nFtSnxlZfiKWP5u7UP+L
w72Io7+ZKQA/3VNSeNVHfTAtwE3HyivGgNx/WGwmBgYtZ6jbwQHxfQ695laPi9Ak
IMiG5moHca4z35NhViBK7+EkLB3x3VrvFZrxb/6sBRovCxhVDujklYJgTYPudvI7
qaAPJKs+grinQjLB324mRjgcfIkJW58knGjMDj+a7QRIpZe0qiGNb+CM7UPxZLxO
0LTua6V7SuUbqexhA4R9VcI2FeXEyLE6O7JrtxBz9VmGvWDyyHxkLCocdWZgHcJC
GrNBLR9AhVVZLneJnSfAQ+0HnHQtGscuhSgHco5wXraqFR9yDsUvsGFJ1aps9coY
xuhRbaJ2oysV14XdqeL2hzS+oqSl5JJuZKwP7iwpueTMNsKS0iWk+LJ1KN7DDcVs
nbPRwtLIesz6zzb1ldFedTOc2g2J/k72ubDKGhkrVJ3/gc3nqU2WB2PEb11QncvN
xNxco1d4gQIxmF4+tWV6N8ug3FwAy3QN45YLPDhwhXe8iM1UbqEQC/fmA/DleUai
H7k+erAYum35YvwTXQZ74p0Fb7GDSPdoNY0FTYIsLkUircVvk9zxWK65q9KcE36O
/bbIu4z6m5RRn34sK0dNsyasg+C41KO0PhaOpgr/gnpB8NmteQIGD2tD3/Wd/hiW
QkCy9HiFmOsYPPrR6IG80ce6rWcWaj759fWPc4pBcbgFoIy3UsbvFO1G6Sw9MfNz
RmsYBXyAOy9VXWIoCIriRerizHyvBtXdf9yNQAjO4anMNxYPZ5kOR1mt8wgoty7z
04//E3FH5S3ZUYB+8CmlPl6D04LpVZn+fbQAp9nYBTKXz5Wm3zJo0ptNRESqsYYU
fsohSpUug+wQeSnbnJ4wELnzDLZRffnR/WjPKGHSenoz0BStGfqZUfmsPxmVkqH4
AZoTdFpARIkRTvJ2vMc0pn8oGoFJfdnBCxXZRuwMoSS+GPzeaWkejWuP/pH27jGE
Z0o8krwib8pCyslxq7wrzmCBK+2ga0zIgpmUMkdzMQAQ7Z3O9XvIEy2/qA9BiFg+
LieSOH/S62+mHpjN/+IEPgtxevhWgcEQWdd6sAjvb3Nfz2+IXAOstdRzHNxdlp0E
bUMiYQeHLHxf95N4Rgx9DGRZ2xudFJDQN/z7wcYkK/3aYOeKyJp9SHVX/PhLCjTJ
96Q9/GFXKtgq54wQnFuFQufYXZj85LRobYVUvpGZiBvPskDLhLzk9/gTi9sdFG+1
pVhDc1yzTYlwDADmepSDNbxZOyTCutfLYbR0mYyu6KmzaJqZ0aDkMnM1Kdh8v039
Gj3kA4dnoJOrQrxLIH+H5DfiBoIFQlhzWVXvZ4hVDf0rxS87pr7FaHbZZaofEavU
rO74CRZofqoeoUChvufv2kLErhPx3k9WR8qBXnHrwXjzYWytlOwhmjHp5yvQ44ur
PGOX7T5+O6GicDLC8+4tDi0+OVJAZfn1oT1FCyGwSGX3Bp7wg9wN84+OFjYZmPHo
5/abuZxx3zSlnywt1iMvMJs7F1NopHUld8K/zjrGTw2I8+xZFFN9IVHqUTeLO/IP
IEsPx3AZvGjCwbbZD6I51m67xs5u0OvfePBZgPfa2Ypnz4jwYGE28+1D+5WX0gEU
cEBxNvHayR4YwTDGiPYy48Od3qCprGqgPyOE6CsDmOLJd9K6/6Y2BuEaF7ig59jM
vKMlB4omIP6agPCmFsSD6L/Bu+CR9GzAiulSUz9ed/W0SM6GoTB5Yq+Ex5RIDHUR
W5fi4XvSvxMh9umkXCjsM+k/YzepH7ENLYJF2Oxi/CleJ2614bt0NDG3S6D2Eh31
wO5DW18GMP1vDhM79dRusoWTf5SVqsX+1WxIxx2UucoFitLZjkKpbuMSqMSEafS4
GLrd4OQuAXLNta8tpTld5pqvXt2J9L15dWzcx7sGtSfsh42DyhTADDChFWeJIbaV
a3yyPKOvxDVt3uT7w7mVSDfCRjnNwJNw4mh/dx1eDy7Y366mJg3uCCYDLFl+ZK5g
4oLdMxhkGqhVZaEvoHVcMLjoQpN2HoveFrsdhiacq3JVueauuGag/WpvQs5CJc6l
csTtmfkD75afMIDMtCBTFOd5tMfd2qhnvQ0wm5t6jqOoOC8sM5Vy5yG4OzR0sNP4
TWebs8PFHFHr6k6whDySDeb7IKa5HgmMsQu73RlgPqCN3vgTjeYkDQ+HPLo6uXZT
1XuMrSAhdnSUO06mipvsD6CZdlayYWEHvWktGy36oO468NedXo9QJe1jWPZfBPrF
H9hxwuIwmxa1Odu2Odny8L5Y1FbZ6UNSe83bSFuLB97p8c9ugALyiblM8rZAealM
6eR1Zu7c46zZdVO0tdwl9js1C+gIE5dVn3zfsPmkG3tO/9XaDUwN3L6Ylt5fu3sm
9CAHbusaxNLBBKAqBa1nG095nEV8rKa3iQD71e0JbQCg+DquaAYxVo+obbOJpQFf
N2QkfrK3aXsdEeQufBrZYeesg3rTbIbmfj5sbhdzYOp7xj+XvEu+BXx1WBAwfUn8
dUD5S/dDHbd8QJ8D2ZbFqmGh4+avqERCRv0COqMs6ZWR49ML5VIIQR27rSq69K/v
jypvhBbmDlxBRqGMGz3G9m4Z0H5gaZLU3XTKq5F28Ye6tthHVjZ/PnHq/SeAGIgz
sIRgKfWRBjPqDp11ksqEIjKiV8YJdRoFFM8pDB5+DU5TY/kz5i6Bbrszpkts2Gd1
w6sByYW+qYLTHk71HaMV2f7WB+f476Dio3Euz4/zrkpCv2FkOUqFxgOAxMmC4q6x
64ysd4ioZGo+TPC5diOoji6NvdxSJjXY7l/K5x9BLDa78yUDS40WmbBrGReBT2fP
RvL2CdXSFTs9LKcW+zDzhKBmiMNm/58vCeMzwDjAv1mS10tYWR8qOJdDaBpy9GRw
IUJqZTF48DUwZY8fp4f9m7XlBVtVgDPxKgkRd1uvcCZEhv8P0Dm5TVcAAsAgIotG
I0Dg4kB/mvoAEWUdU71uZXEQlbkGe1CwFnYeEdgGgvej2Kf8wFG6zeNtH62lG0Sb
yVzKpwFcmpBsXrUreUVMoczJnZ6DNkGTFVAoNXLgfwI+Jtlv79jCoJaOR6i/VCv0
cPXXsekdjTut4aEHw4t+Wpu3sjhj28FqGupnzsX7cou9TZEn2BvtvEmCsbNOakyP
8SoDVlukY5v9gnDchL/ipBCufRZRS70NJ9btAC383YkVOZxMcmvrAQhDtdm1Pt75
DZCEGR5skwrFB6JWv6f+D+CfO0DaHN1waKaECufy6A3xKFNwKr87xcsfHFZqSls0
0daRYdvNh87uRRperizQ229WXvGWU8sq9RI/as/7zJoltLb4JJn3RwoTTonyzVLu
U4BOECfw7QwQ16pclnmkZyNbt1cVOy3lLV82npQ2rGkkTESvV4dGgqn4smv6Ldqr
/hR7L/dDrPHPty9SRH88hnjhU+Ft7FL7uf1QVdgyYKD369BFbiU4m7ECamz+VqVQ
/Eg3+N0p66YHl/HxUlhetVTaOTf8IuFEJPqL2UY+cQ7CiMJiTpsrUhgQEVxIGUWB
fkTTaZU/phHWidgeGgfNPbbaso86ILBXQgVdMG28rK4xqLjqtqDae868IcsyAGEv
XZKwmIoj5dipHfeZzynCf7H4jx8CINEiGz6Kyl5vt+SwyxGQJO46Ec8WhhIlJ0Ln
kuCOhsvL13ydkLTVTXdRYm2RtXeuz5qxJM+O9UVrHyNjjA32fd9FFGsE0gpdvuu6
8o//o1TPp3hbeNUjiU8h5FBjn22aO62ZgBkHUOtHo8YXnKXZPlYRl6lKq37iUg8D
Q+AIKKHrcrerDzgehGEgUN+MpMbnu2o0DTekEk7JhM1NdugY/FcXT8fAMPklDaBD
B1re3lMSPxFrE57NF+5+0YW5Vpclzd0magkMNco2gTFqwfxDD0oopUzGLQnINyU8
pm+NvvSrI+Hwdvzq2tsc2r50ry57jPO/XhZ28O+DmEM4XwTypTTqHlVI1WM9OajU
MuVXIrBTLN5FGbpB7wuh73yz9oad4lEBFJMqB+bVkPPUVfA9F51y9G7UZE8WhfJJ
rV/6HzUg1U6a8BOw4+LAZWKOfTt7hw4Yxyx4NLIqYzvSZVK/kCc8OwkqfWCAJFYW
qCMstl5PZWh+8HD/fle11FzNgWMFxIlEEL8OiLcBeb0/DhhZfTHiZlG+WH/U6fvJ
lu+TJLDnNoRe3bguJSWf1DYBBXfp2JansSVXbUvObYck900idaU0tlms46NeMhjY
bZv1R8LpJeBLHq3zHypxQzpNY41p1Y6HnwZR8NznZZPdOUPHtCCKd2whkWEckTL6
ke17TvlUgkCmgVnBH44ndrE5MC+onzvCLUf0jYfKR5evYmTZzm/Wf2NN2eMdmOla
SCqVpIfXBw3S6bOx/CWs/2httz1ayIB/11FIo8op/IujPkjcLlJ7GB18ePAB/JPM
Qx2YQo1zzJZ4JDDnzokuZafxlgwiA7i35wt9bqiH7LP0+ccXEiruG+kGrkh+HkQk
VJN/8/JfhsNNEk//lu1HjEySht+TZ+72VUejUJ8nWs99u+ZjFn4zrZfjctO7YBG/
SEzfywM0t+OWRCwU/DRnKm9JrDcJrANo3Xi/AkVELWwxq5kmr6i5k20yJiZjpoET
lQJOoi+o4ksqTXalkmRCx71rgMfeiPWbI0PL1JAhrgjzq/rXcBgI0VgWKKdRzLXS
R+KlvNKgouDkbJL7m2hZPiAvp4WjsV0ywEGgmbiQ1+1rsYjxydDopjhBj0M0Hm9z
82mpqi2SkkK1EKRGgsFWKeymey95RReQltBvtw0eIl5cVn5lun98iGb1EN8xB6c0
G9t0LU5GbgJWL4hc9xfT6KNmr5YhAiFXiG4Jd9RIzcs6VjipRbg+1pgx8OBHmMd7
Bg3LeovOJv18LqihFc8zPLVfhybBIGkn5LS1xWPFvsOkXq2P6ITHkvM8kqbBBaTd
2jRtTgCKtEMVVAqPGiE08dNC44jWtoWi/mV2c++Y1WrMJzxYHK65XF02dz020s2+
8dTjrQcJCoDHVL2Dbek28ISCzQHTCU5SeT/piKKAE6mZ4Jwfk7LTA4z1aiVPpkMw
LhiQpgQF8Banaw3nMxbdBeNrsJd5SIKXNe/wQDUWOkOBTleXx5bNAQ1L5mTpFP5P
G3RP8yHMp8El9QPuV2mvwlmPU3Dd9YwOhFqyYgGmu/HOvcPBcbQ9N8uaZstTI58A
gG8itu3U+yzruTveAqSlfq5wUqD0qI8QZyny0wJBEa8pYOIgQx9Ltn91ODVTkUB9
4zzVcYtCX1LPR1/VmvKxu0l42Bxo7gc1qRj/xEOS1uVcfbSv2MAYRc94fXGo8Olw
CsmH5NTaU8ixEyUa9DsFs6RWmVd+PYEzerz6meee5bOlX4K1hPdunR2jR1hVouZz
qZE2qMXGm8gFz1FgvpRvVM8teODxipman8ookPLZ9hQ4PbEC0j68Is+hfQtWF1aC
YCCe6KM2VUvZbrrAl+s3rh4RO28/lCWHOwVjXGQbtROc0KYOSLe6gL8xoWcnPAqH
XnXsP5758tOXbHWB3t06DKhhQId3FtaYA4iprCz+k5oI3xjuJalkwYHQPWpebAOf
0nCptRhKj6md3iyPR0K93Aklj5ohQbmdGOTm0X2mFWc+nPnzyDhijVf8RXbC/dyD
rBePj6ZhosR3vmLccMHxWq5uwNmevLSDQqZlFXmOaw4LVTwFyXVXDULOPkm1g+aN
R2lu8QJgVleqIZj4VaF2L6Pfa6Xvmx4dn0YvQ1opaNDqcg9tEKJ4QOTZa1XzaVYX
Sy+b5SX+MKwewQs3FKu+SbRXXmiCyuZvJl+CspmnI/O44FozxP6ZSsR+DGdBCQoz
p4T/sBNNW+jNfouQ50GnDvyrQvehMWy0tVAAQIMYNG64rl+QxWixW4qy8GdriIZp
UKWzDNgGLlmcF9kW3iLIArACZ3uVIUvp9fYn1OC806S8XmyQn2XCIeXOoxOCwzhR
Te0fd35WvIfBGgjOFO/3eO3xE+WmTR26JiiQdapY8CRhnDi5oJX9NnFFM3+bWCax
GaLPLGKNT0nJy3a/aJOkWnimXPcc+N7ZNcVezYFS5e3jgCSfq1DZymOG7bnMQpFR
3jNsUVVSNWIHizApWzSry1A/dqQP/bnUtR5eiiIryd6AiqD0pwEqzEELgadN5y6F
lT3Xpwwap+3nGKWkRPvk6cXUhNb1xk4GSRTJXOGxKxELkhPklf6v6mMk+Pk0d5Ch
xYC913XxY/2Vi4acIzVVrM4BGLV1T6ozjbSWXuGq8lsk5w6/Uo/Vf/PkpNqy6KZy
vgS+Rv0XSia5j9o+oAhEKmj6Vj7kaSyLYV+mtarbkTCGoUp/YGnbcKvEx2qNuwCz
N4ZMr4T1mQHFQxZ8GsMUdJq1jKrJVircII3xiy8MU7EfKinlX5YALc+28sayB/nQ
p6wn5wq2hYYU1OBy6p8HRpTIDgpaH6AKoTSEPU9Whx6fV+WrBpaYmPHxxsq8v3gW
XxF9bk+NxSgR2CkGe4Nt1aKXGUwo1IGzIyrBYyTA00+0laSmjrBevC02UTN/cbTE
ikanCWJeOhb4hfhxYXsX6yOkBFE3KzIKUOL/JMxpkC/Nff8oyldSIp7JwkhErcWz
HDoMKrd/qc4UkAZ6JVoRkqSyACb0laz1tZnQOoLXGjeI28Rm8UAcmFyzBlj9wG3z
F7+Maf24xhU6x9SniMdELarpbWbEH0mbsm5LLHPbUVllj1LSlBKoR8eYRDEafiEJ
WMRWIZERtPVThJICZp/lGBNO1rBShhYtUohajkI/yA0S13vbYuCw9ZZETewhtzd2
VPE8c53zsTpob4n/nnzZ5TnMl96wTxQLeTKP7/USlZJbDixHk12IHsYZ+XpONfIO
B7oc3BspAX6AHKGpBpBISQk8oPIaSOIQ0XO8AkQE7JD7m7FHkhpjIjyx7Ok57UCJ
3kMpBBLtgXRCWvn53n5o8lQ0j9kccHTrA7H7C3zzwrWgyGm6N8eYwo8/Cfbo+FE9
DG8W3Vl3+/mkqsgiRnHmZgGF99LA2zCagTnjC7TmwaWHQ4BwfAAIsRV7Hkq8Wfam
7zxNpwD4LIXncme7aBbiRsKGJZXaDAm2WxS8ffdqXVj84Cvv2kEwrD0PA8a0kICp
uCfI4/E7G3Pg1pfUzlvcJ03nCoGKcXyA4aDgJBYRJ+Jan2blabUn1gqtcagok4DE
p5LIWBv11QNkx1zsaxQx8glHGx/J7rSHjRA+ekcl5rIeNh+fZ0g93VFx75tu+B5x
JA4dUgPI8CT1HKwK9YrQygryLZfKwEHzXMpbFUBHfhPeYuZlw4QkgpB3/oCKeqHw
GzCEqgcjHkxgdQb3TWdTaQfSPhzcafHM88v33pQLUq4Butve7LDvFzxtOtBFgG/f
BR7xTX+loVIV9pfICMZq/jPbB4MuffxAElBO4cHQvbVBjO8pN6OCPsjSF+d7e+Ly
WkPQ4vwyzW2RM6256SHJZO7i+vhOYmpOdblCelFL71bGFy48vAmTTaCwTssN9Xtt
uNUX6RXkTMM0TZItItCJ7keAXZN2zKEEysb0jlIyBRP+6PyCd5l1bFxVqTA7al8u
kVVAy4uWST7ooi/D1OduqK+2We5c/tSdJ/HawwcrPygnYVBfLB3nP0mYg1Xo/mO9
H0365QPIzvPMtczp4LI2Y9uj81biJVA2pJsNWyMfE/Ev93F8K0X0ljJz0XHsLrxy
rqbJg2FDCwo7B2yLQQbkkB3nH/S+3reEah7dcrrt18nRYjbFjIanotcUgeyI6ZJ8
GMk8tM72J43kdMasJ2TMZv/NHU1YKQYZB+pQODdOEbzUrFUCUDc41SSSP4ArA7Cv
FOZSDD5lRIYlMn3x7yRlbsJA8dAjOU9gEu+olwaK9twn5PtxHP/wyGYAfElD23L4
DFSQ5EEpSs5pVwOqkRfX2HGQqRUz7zgj/BsxWbiHtD+s4Y1qd05bEbRnJX4Jatmc
JMnXJy2fhk2VvGWCw6fv5Zr2l0kBCHzVaxDzKHk/KYirPLSVmPvhISOhHng6ixUC
E/fQdwgPH9vHjco1gxdyztWlSA4FXfYwhFDXI7Y3creTXx5pBH2GH9eNUKr83Zdh
8jWTPnIEllxffXxbz5jIs91qO5IJ09Rh3bxCBD3EjbkWHtNVfnUf6Qx1P5MaYn8X
5rfk+2W82F+ugQ0hgWesGXeVjkVs99ll/N3RojWVqaIssa8y7A+f9fODjz5FKRob
9Fk1ShbW4oPp1dQXCJnDP12zjjRLTvpLsMKYAFQoHltLI381niUaTOd0dqEQVYC6
y3wxCkwJhYjm3i6Sk4wAaBZvZRQLz+oM8EFwiQaPo52l4hG9UE6fRR8akpyVigr3
40Z0gk08344Y3Ud6YYUIlwyZcXsShp+HHJXi8Y0RRwrJ7WmjgzfECVSO2/4wqfWJ
rHx3vUQPClayIG7l5nArSkVoEgvWTSmVsVX4NAd/LFLIEmU9fdISc7VfaTa2hdjb
3BG129O11HVhMA8zhp8ZH6d+4+52zwnHjbG4U5Rn7f+AylnLgkR97wmN4cBF74hJ
h4r0uwJ7EdQHGY4XFsJ50D9JQcsaL3OUUY1FOOGLsjjhRzPL5aoQjmotDMChA6YU
qPPfrkaXaf7zOgX8aPXU+EbZZIgqrnEbIK4whBgE03bhLv9ucmA8LsMGPVj/vG5v
d8pmW/ACJzP1BAygCLchT45Y7xrY5VqhBynhtiIWV1H3tNtuS8eTV0R9zl0bzQAm
E1ZLd0eVWkOrRPU2Mbr0jyI3Ec5aHuQirH1USiFMum6FQK3PZGg7as4U2kZCQaEX
z94ys/akUYW0pDtvdc5tcNVZB96WyCA/zTz0NK0n1EG0Gs+98gSCmifn/6r6fC2C
QxDGQAG2XSMJrbijVhZHyAjssnihlZNfHAeTr7BGwRsdYNYv33RhqhfNZEQBLHrx
7APZqdIQQurAQO/0df8WLmbCFqmgtOHQtZclpMBVBBTk9X7ryJ2o92uRssjSVDx9
rvq0HsGW1VHutf2PzlNHCa/M76Qlvxf8FuFVgC3eo2KJ5ZqcdTU20D2ahdSJYtBb
acVSAGLidg55FAQBJgO06qB0lQ4mxoM2k48HBq77TPfZX5hHvRO+/v3CHNOn4hXx
Y1qnftwDdF9YoVrHtoVxW+27EVc2czJvfm6YbxzC1dZfiHMU58QzhOXtoLYzQm+j
YkbMKHwyc7IPu0UFpYowJHTxtoETELnFj2awo4vcuj35JfQ4+npdbyuxggj3yfTz
hWabqxLqVisohdBXLn0f6Eg4wPBNVaqjSANPP+Oxaf6i5sVwL7oxhxZVjQkBaWGC
unfg8PewiVxKnuKIuoeP9QKPjtR46tbFxcjczZ4TaVT+62Hz4kQgtDgEyTSeIW6C
42sLx0rJAWkvcPCavjcYVcdwCvhJjywBQbJg+kwXMtCe9xIzfeyBrkZf3Gk0d78n
uy/G2HZJB0HgCoa7UNfYd8eMLsbZNc6pXsOv8OkchCDhIDOuIKHnPqayyROT/jjC
97SiBlMktT3JUEblbsQ3lvOzW/bEHqbyhFsNOazp//W6XiGVKEIp6N6yL+KYXXKO
X3VZ4usnpi48dLPstdbagLy9Ur6rItIHeChBGJM9pc8GC78mJzgYvPPowXQK8F3r
XQiHz9ljOxuPPrQuUB4TrChc2559GU9/b1W2Ufsf/u5ozFSaxSNwcdSVZQM/Njmw
gzDB1zNAE3bDZbNdzM5vKlUFj+MlDPgm3TMlnZ4Z25qkO6pw8oxS2b9PDKb/6yaI
59H+ky9MPCWCLfbvy4HCXfAucl63SXDDDYPDAeJ3zC+VXY83kw6PhUIICiA2VF6X
3a+MuRpudtIK4fRCS5pGcPA4BwQeYEew34H4dBTwCm5vrp0oC3IKAwKN1Hp69BtB
NbY8W0yO+IXi7zYsCgTUZKytOYrNrpgh2m5IAUGcBs8ShYn2mtlBGLYmuSFnsSuz
arYKgt2Nc7RutAeEQTvN/DEqtHtV2YkY19ilGi+wVTIa7CpxHbUDC1gf20AnKple
bnCDIxyv8kMcUQnx6OW/7NViioPTsyV4fuCv0Smwtc4B+e1nkdK4Psh1NwbpPZ5L
cc4Iu6dnhOx6IZqGql4gp7CRajsdMfgTBs+usY0JOjcjzr9RdS36ynPtIeAtbASL
WGXQVeG+pfPp9ctUBufhzUAv8oqLGIePMcd6Hk0uwIdkxvz073TAJLen70H7mnqx
9hc8bAO7Atimtw1n6ksXlQdR0KAB4aa+x4SBoL7kut8/JmbVdFh9mkj7hDqS96YZ
+JhEbTgXKN6hHOqLzYx1iwd1daumBpavF0m/LXR9QpvPiAjmv8KYd0qPUMp/VBs8
emVqn7XG6qbwfeZJKdb19z7klkwNiNKoWrqW/8Vz+c4jda1eQC3cJ8H1ksMOA4rm
nxaMzZz7/ZmRG7TCAZpmbu+JWyTKkbNgbIKjYh4a8uwYi8i8ZwiwNcKjxjK25Agz
pKArxJux3luG72MrmGjaHuR+OqAD779EJn6pROze8hD7enr9UMEgqlZdsmDJP/41
c+/HnA592JpWSW8NIQJk3QePlJ3YytxyPnZFJ0r51KwU+rB80UJXpFwsqauH2E7Z
81kB8ZnGx7MgETyYXeVfuen0yyp5eRn0NtCsjM8ZOGROdcqCPTFx+zQ1hP/TzDAb
MIwwXZ8VSHIpJWlgoJPbAmFH4v14vw3P8hCQd4BhOfy3T5dDYgYhUjUvuwtwAD7/
SsMWk1CR+mm4fs2JxFmao9XDZkD4wD+1XTxzwkdcbQdIm6p1P8OElvEySB6nQwOb
Qw4EcoK3WWgkE5pt20n9m9y8nanhKRfmjec//4xUap0AzLEx+hPuTtx3+UIXv+pb
3mwCh5+neos1sncBWP0MFz4cVYiHfAjV0nfRGA5xDr641UM3hUi6ckaAXGGR8EzY
WUMXeGGLnNCJgq8Q1bzj+A==
`protect END_PROTECTED
