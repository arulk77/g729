`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFXGeZWXSp3XdY6vlFAWw/vCWRuKwBzBjj9phYrWsXEG
Clncl0ZVa07idJc9ODybiuBT/CeNqhelBt4xk/jEBBFvKEV/m4xA0Q77XuUN6Qdh
yNxZ8NanPh4tdF9+Z2ihWXAe5wysAfT3OLkIrEi23ZypJYHEXBtEDf4C3B8g2gBG
a6jUyGco692DeX2w+ge70YfdPWiHpwiWgbhCBtT+3xzeIt/HOUuV6HfWKQNMoF0n
xWkWJbGkVVpwvFh+dku+aDiEB7zgh1YUsiP2swoV4qYErb+KEyx3wJRdezqoRf1p
5gvivxqCNjQBByfhZaNaT3cltDBcbq7TG3noOT6GFiQFy9pJYlZcRqOs6crx3TdF
24Bo5G6Ks6irTPr06DyAwMjV5x59aVCTvTFrqN43dPyIp9wolVSkQiIluNRkc2gH
7KnFOlLbE6+uDWh8swalStAkq21rbMiJKn1Y3a4tHXEN06HSTb/Mdvms3cJZJcE7
HnnbXS4quWay49eVnx1cIQQX+PRdL5ZGfWIK5szGGTZku7Cm7+QP/SmvI8J87L45
KxWUgTaMKe4toa6yaHyhTKCvZWVYG7Jpoz4ob6VcY/Q=
`protect END_PROTECTED
