`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMbekDMHnAhitZ6r0wJbPKIDQmfU2P3J4GTXRSms6nWx
uIPOK02Dze9fcfWNAOcZDuGvYWNLRUSuHmqKdu/CFn179dHc7enWSPVI8yjW8HU3
c3FX1c2fBC8puqxxwoZJBztlBc0RXLgvYIpyYy1oTv/Idud3eSkYA2uefKOgUbm4
FYFudKCl+aXoRKcpiLfgNw==
`protect END_PROTECTED
