`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43BQr61lKbOzb6302gP+x41FKnJwwg95TOf7reHOx4EU
+aI1NZMal3ujBBFDeb+Tcxya5MyqhvF7SXWzfRbUTvl+K4F83T0MEmiptKe+lpQv
wqYeuRy3Wf8BfH2SuzDkMsMBggAEarwe4p10yKvLd7GCgt3xHiHo57xxHl+bRsZc
MgmwiPlr0n0WN5PottUs5LE8fhxnp2Fg3ZvjxATdp2ZwrlTyvUu4RheunxOR5quO
PdnE47MO4+zDaoVS17b6a7jqi95IXBcPBZGihx87eHsJy35B5m56r0OiGDrl/Kmi
eeEuCkGzeYLJCQzLidR8UtBRsbPcOTC9m43nqgb5AmAOHPx1zGSRwTgYjVPM+Qsi
nXzBty/3UUuS/FTWvWIoAA==
`protect END_PROTECTED
