`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN295WwdTxAcnWR/LC6vb+mPG+VHA2o2fZD/t1U4RvZJg
AReZjjdBYy/b3Z02mQrg5oaygIDOIwcKse4c1vTJdMjHa5c14Xeh+sfhSueFqbCp
aYIN+mArBU9IqmAsrCr3ZQXqyNdNyAo430y3Mm7mhCrzaRXS0NfhtnK721ptDkRu
/rek/hoVobyjJioSBq4OCzra/BLvD7v5QBUoU7YxhDIO85OGO8x9GowOS+Ah/CTy
EqW7BHVcjEZVII4IcpEFI2PHECtreQ68UKbTdaZSnDA8x+GEIGxtAMstJ+ub++dk
BXEQWi2VTVdKWCLs5zYQIddEJAsH3GWoldp0mzZOdUBoqAYxeWzDT9Gt8BiVkwHI
Sw1AmkdxfmboBXP2HQwZ2n1sI/lSTZlb7sBpxSAZfrrPyLYePBS1mjDaw4x6f/SG
FmnEzxer+k+b0LiDaaZitD3fIOraAUd6ZmfSymcNFoTzyhhGDogxyLJLNN5hOWx5
IjwCcDm3ssKwEIWtMoqnBQ5I140rz60L7/q/Mhyz/I0GHNLxFbJYiuttJs8OKUJ9
0risuqwEhDsyynM9d42Njfj9XcuA3w8QVGrMS8vgt/kYJX/33CLKE9TN4mSK+ctY
SmUiRHE7JtpTSwKT51S9IqUglSTv4l2QbDg4dJlnfu7V/lVSBjoolgk95NwYIWtF
w21Id5yRM5aDCJrKTrQFCOXVsiEDs/jsXkWRJwYi7dRqyIlF8ZYAoCzVXtxOjwm9
7Tf4qw1YsWXQNZC2iG+kHdtKX4zry/SzQk6hwFFScS7lQJoCqEjzMYatRbW/7IGB
i9lhDKzUP2/i0tMdq+d7mMwuU8lOMIqnlMy6MmYhHgvTdKQKLFeVA+B1ijhM1HzI
1JvRTC3e8xOG2izL1jGsZ7pghk1Pl2pKcS8Yb764RDW6fSMhWPt3uMjVXDG+OzY3
+nO6rrmApH2BfdfmC3tYzdlfuZOQLMtPbylBGvLVGlF9f0/Muvrmic+Zf3Wql0wp
Zt0X9wcm8sEr/n3GVsJy2100ILyIk5VsC03Vr5Q/AuUddmaC84orPYp4ar2ptRNb
a15aNTnF+pngo4/zu4RQ4BWZefchvCr02DaYVUYYtX8HxuHm2+mnfPaE0pq9bIit
9v6nMOrgyJD5y6IBlsYbQnsbjgrq+rTc7TkrlhhEd9ysvrIHIF9HriZ1cqgnamm6
qMyz9qfHwOm9Y7lA+S73Rfzbdkwsk1yL+BdQUwJMOQLfyzRaHVa5Bh65UB/2JRsM
M9i+/9B65SgH8nmmGxOttrPNnbwJN9wF03Q1A7QdR336kdQW+MM50jdrGPImxoBq
gLJq0eq+RjuH30++HZ7msZIrtT8ASh+MlVIZRGtKjLXfqT0h7zihfBnSOmXEohFx
qFK1dXd5+D2FZqxoNGAG7/74oQ24uocSxoOP0iw9AArcuN8zwI6zNYSFg7+xgHUB
vMuBgcZ1dOLIlNlad3PAGo2VWAfR1bvWqwpguHFkt2RIHpbayqMHTFeisCA+n6ws
QIxhUvQJ7G6+1d8nt6IfwKIk/rx+PG1ltv+RScOcg06kpfBkGpUCqgWR9lV4J2up
cg067fXJyihO6tU35sStPrwf7ZLK4rWsxqag7OoWxItRuo861mmcZQeBdJAeyaco
sc40S+cMS6T6HY6xr9/BDq61IsFA4Pn5Pw5rlrsF8e2XPe2AdhMqmh7fe/opzSOh
PCL2GWDJCQfZXczS39fkNkjcGbKXXXmpa0ZfTjYHhnME25BClFePRPt0OImxRKUK
+If4FjIV2vtQnqRApYk98fzuuzSwgoUaN4NKSMh56/3mvYwOGi04VgBcMEeWfiig
GOiTiBgjLAU6kdZjX/jTlDj/oDFMVVFygr0FxzHa2EZJ32vQxgykPvOx4A5O+Hsh
vfIrXnIhysog3gh+JzIVAQeVQcbVA+udUSddtYZwNxMDpZizfFQp2sPOKTXQ5+ci
spD/OZ4BpLhZUMTPW+g40hh9bTqqQfDJVMPD4Msw7MHnIe4grduXVg+ApLTFNOG5
Z3BVcNvJQgHX15b6evYyMoxTZlEtPSzWOT2xQNJTLK6Ckc4B/rDl5GUS8nkwooNe
y0B/ONkXi8KQoR9uH5F0fYVAGppDM4PGyPJm6YQdtx1PPF5dSEK4eEaZLBTjnwI1
1fPPRzCq4pJK/a6f2qJ43CsVkj1DyX74RaeJIkHryzGU1I9RCnu4pvAXNQp4b9wc
6qIPdW8lg4lta6OvAaeBifBv42XqpgRUtEWL67jIyZfuIY1i7VQAisCnpjfKeY8I
HIarkCXnS5gJGczqe9nJ+tTnnO/sPR8axp1aTbubCT0099hUqq92TIQ2gg8izBrY
yQLVnOhGJcEoMI9ioBlQrRxsTB4KnbbWfpNTwb6tEo0=
`protect END_PROTECTED
