`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAcz/XPWZ/a8S30rQNBLRzSGJRsIXx3u+R4uqns6Lnao6
2uHB/GADBJyMbVdymC/88ka/01/9jM/CkmHA3/xv2jPDZzh6Y/3MBRTG97KdJJnq
m5Y6G4VsaLlARidbIB+EF7kDaozH6/51kxRQrDE3OC+m7nud8jfZmv49amO0uLVS
Z24ZB6epg96ox4Fi3F2WCw0cVE27TG++VmtDNorLuOHFDDxuH/Wx9mqDhVvzGnDp
V2bkgIqF8hpPnGmCdXAeLdK5jlpLwOzFnCCZFtM9M58kACLBYoS+W//jUeo5hpCM
uOpWzlb0OGf60sn+81+6kFgiFgLJvhWoHVF4mmEmXtk8WlesQeG0yO0ouXCta5+m
nHGIz7zjRuqaMjNmNfJMinQb54GNtgunWyH1rvOo9xntTGlgyMi1Fk3/ZWQs9LvE
M9Yl9lDL8xD8aU6f2iVrWh5HlE0OvTanefZVSYn8ww6og84jVIHaFIxHwtI7BqNK
GXfDx7D3fxAOxubZ18TuvTCYRFQ4x2bqqZd5fA6Dumc/O6EiGQxq2R/JnJisrl1n
2GAiYzgCA6/sEogGCY+BWgc5szqSxPWVcGTXfIsQkvBC8dmKQx+HIWprJntT3RwH
XeyD0CUya6gyyVlZDbaFEifH5ptxfxkhrcgDVH5gteOTRu6H8LD5wXDlJ1kZpeLx
wjHFzBzF5oVp0UrBc6Nmqb+rfqOXEY3BJbrutFdDeBc03jWLrtlAoF/kSLvx+GXq
NRWTQAxkPpn39H8xtAa14SyG6hsJgs5YmzatSRbrARx3hARWiQ5M7d55AYYTUGNz
tRkHut72huWkoHb9BsWLCKkX0rxM1oZd50j5WOlA0aQryV0q9iPYr7uXPWsGtCM0
1lvYQXDcUd6D9W+TKSayCBWEppnurGSh6Xa1FbP4UY8wHDKu1gwI5zAtKo81wR0k
nesJ9c3Jwd6qnf4GYmmB7tu/zGIfxaC/G3/ZvpmKNmeupTokny7fZLf38q/o/prh
fpqF3ZOb1AxMA7uzihkhqGCPoAB71d9qC2S7CxrK7umI92xp1FM5aX2JFTPuOl0A
ATvkXbZ86MrGO4X7Rxq+hmNSP2l0SfyHmjB7NJTNR0TXPoCXJpH0EbCLTkBfi/T8
oi/L9k7PQ18KTyGoRYovnIe04zbYsdOpC7/SWsUBPvp+JgSkpF5hF/HmarXdjNof
jQS9nDf+ghp4nQp0uTMuUHlw5CFjfVabgYfn5VkHygyyMX/MhyCTFg1KUIqzdSAE
Ipe8jTOWfNLZu+yXYPhVybuajAovoi3Cw3J16Myw1r1Ie65KDXN8novJq9kfai8+
erFnC9bMznllJNEPH93XhYRwwiFSKbXhqaQl2ieczSKj611Dx2NOI28zfW6KUlN/
vNutCvJPPd9sda+4r9E/rLnlRlM11UmOt4CO+x4nftPt+5TTmUpcNGZE7e2sEwB5
AFU+ZZ90J1Cfwujc+P6FIET43wQfIvw/oZJE5DQcA35dq/J7fxbmSAxlQ29IEh2E
Q1HBd4zjZL72CAz7XwXIAzHkKdWGdgCjMc8WEPHPlZxMQTtZUDBqQfROAx8zUIdd
iAx6idmtdkKs3taQ3HI4uYa495qp1Pn0zjkTfMOmo2LEIaPTLEzejtBt8grDmNsI
sQUOSUQsTr59q2XCiV4ymB/bV4P7S2HwldaW1Tjin4oAy/rBSq5LgdXcJ7Pou993
nVBIpzb4pvIHooHbN81ENs74wih1d0Y24q4RZrS3eUn2ue2sjmLbt84p4MguBdu0
fZc/qs4D9kKCihekooBiHgfwJgrS08u1fefUrdQaHBsgRUNeY3/WILr55Haa2H0s
VHTvL5yLkgqs4RlO9uQ5RCEwH/o7FP4d+PSxtgieSHZHIqzKotSRPCmDp/Y3HEeD
3J+im3eTRz5cO8Tf3n8vCRMbBVWi4Ja9LvjsbzSJ7vELtxXmT6Eg47IlGCKxt62e
lKKM2q6pUpTZUyJ4mOOYj2sHNWxE+gHM6EqunTLUwZE8L3H4oRF8dNnls3iMGFfb
YQHTCKw8SNybzjsVGensjywvhWOXnk3Ku7tflDanagUWneUqTIjCgR+mnqRsOTkp
pFWTdxNhZ4GTsYK4AUG0WDXlLgfCByT/eFpc0uV+NYg25Pb5GcJn7W3P97L8XZ1+
QBZuUtoVIlZqO6KDj9MC7+p0/BLvOYZaAd6SlXz5gDS/JAsb69ogVvw6O7oCcPrr
I0b4euIGkq+Ta/zJ7Y+0NZJ23RoKnTnUoFPJ+2uKmRbLcUzstgU2gZcSikYt8Cri
5w0C9tXcXHQK99wkiX4sD+ZomPcTBq5j387mMloz1BtLnorn4X9cDgH/NjvsB/b/
oIx/si+JzG20IbucSM0O5lTatB0e0knJVrYnfflRaZ1IPpqUPjPX0E1sfVri2ztO
iurywbZNBb7zEX0sg5NhJLIQse67Pj0iljp1dEXyBLiVYs5yPjvw62C7Jbd3Pmz0
nOq3jgoIJDBRihgneV33zguy55XQ55aln0bAh1dhnYkZDmLKvglwGci5jeAIeiE6
MuGgrbqnJzXm8RRlS/gLhotgkCKwE6jYz9vySA9/rTlSEiaq4M+/GC9yY00afa0R
0ZmHlnwTePkaSAXfrzamScn5lGGQrtfhPixTqmZYMjRHBsRLNmtrrJOuhSC5Dk+P
qXUuVuPq9W3QsPg6SmOVrzfwvArYhu4xaiIT99/XipbAR4vX0j23NrKRlSkKOAq3
kgF4fKLuE9c+TBKpPWCfJqtw5slA2UacEKEDjes+x0ByoKdCUHXJJDCsfQyYyepd
`protect END_PROTECTED
