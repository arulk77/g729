`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOgGkn9Xe/5/25/rAbco2orwJonS8x4q/WjDw3npTwF/
hSI+rY22o3T2SRGPQw76BTfawgSv/b76o3cCvVz5dvH+b7n/AL9V2beYIwDpOHSF
19Aos6MOCyDtPy35mox2sYD1JOyLki6uV8+l7FaS4ZFBEDaJDPw4SbXViOGDgM/A
FIKxDSdzdLDz/rvh4YMc0GsQtRumppZ/4nFxC0tuV2IEyqvKj6zZlw2g00HS4u7V
We5BKNz/V1RpTu6P5cnGQDM0vikJTpapmYG4g9qbJ57ZU2ofISPygxBriCZoNNuv
LZRc0D1End+FR/JyYsV3FHH4ADv9bS66NsB3xNg6/VTzSZEbz2TA89kyrJxh8qYA
S42libtKGjNvCWSOdKlRcsDPXcdO4K/Q6iG8pxZ3uAtEkJdabfvrYJxQ4cRuJ+zD
0jnNox9YFalkQW8QcmsNwt5QzME+NTMz6xo+GRlsFK/ragpYMDP+/PByDjexHJ4z
np38IuFuGCS4I3KwOybj/yqjZsp5SGKr2RUu0Esxw/E10tWLUx8NBxwP8TIjsQXn
24aJE6eF1BKx+ikl62m7gIHe5dkitSAU8nojQQUn/mONXV/QWzXgINHCusDr1dKZ
Bo+WfTGKS0MPtFaeCd/JC8WLAoUqAZPfKjP58OO8eDtYVDzOvI/d5q4CG6gVwAi2
`protect END_PROTECTED
