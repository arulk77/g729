`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIDudAy8BKjs/ua1HS5eWclZe+kb5xiGFUDy5fqNZAYS
ZUXBf/Cek38Nk57SjKrE310oZtOX1Zn4I5t5VRleFTY+SxcFmqJXfYh5AYzAMZ3+
nEyUpLNpEoe6GT0qMYl724Bh5LkCHLvinilJPPGdNK65cHWlljFRgcHFbodZc3vF
kFIVtdti3XjdI8tZ/01djJpcmLz/iLOUXcdig9DquspDBNX0ntuVbAr6TEsCWLXO
`protect END_PROTECTED
