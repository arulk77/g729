`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNXJu6NB7WamPA0HOb2BF2dl3TaeEnKr4Vdgt867PmuL
VdVBL8bDZ0bka44Dhhd0QsMZyobgKlJ36mQdyHauPC941isPvKNHuEEHD9bV0C3d
wLIV80BjlfYgbvjDNrb0q93a7isJU/9mvgTyVYW5g99eSFDh9L3nq5uH5hGeJmTj
SK9h3kax0E6ICBrL4AtofYm9G9MN2F44b1zXF9OleDuKGVxOR4t7/xk5Ml/9eYVe
7Hn2nxvqXnAxNTxYHIN7elsD/y/GJEWW4FqsOO506OOnOuFq4lqgP10mq4u3guj+
qJ8ea2q0W3x/83ejLZR+3g==
`protect END_PROTECTED
