`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
sLQUco2KscOqI+T+0ELAbBNYGWeBi+TMFqNjcr6w5fq9F9d24yhdzAzhfn0QaqEy
cRmKwmgk/57iKfY+vnz2E116NQ9uLWCJiAYQwjxZJrnWUOvQF/1GEWO4ck0N6Iln
QA0REmFjEUn4tlRL+jn81b74YFsOfZXRYH3LxehRU440+iLfikAgfvBHTriuxRiJ
86Hw785BiGWfYbmHWubc1HrAWcu72AnW5757Gy6Ai5jVqrnBCgAfDVsbQ8RpVdKd
x8c1tzV2tHqEh9j7U5w/8rKdGzVA1vGKV5Lr0w3hvbs=
`protect END_PROTECTED
