`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mxBB79TLPe8DY5dESmuJkqPpTDgzPpWWPV70c9qNLJSKkYAYnMEsDlMvYF0rpOiH
4YK4IT+nuswv6sg80PotuRWmgy9jBwmIJWMXueKQ++nlbpBp7XafqOYbQB670xmH
f9SKDaDwQypg0T6fwnPaOh1ArcHL8m7zBntkiVUJ3OfNN1YHvt3E3igmEbMPaoFl
sdDnxrIUVlBItM4U/8+90frd/cdcy4uJlSEuyr/9i8IkJP71fcjlX1+X8IwfPUO5
tqp/ox2KxIapzZNi1Jzcg1Hsm/utgSSdzJEVOC20isU+FxasPhC/F3btK+Fz+w+q
3FuGk6vKHz/gwpf8VZ8dxnlb7pMfoLS6JFSL7pGsmTNTVp5wEmeShbfr30/ZxMpU
ZjSyhxxy0xR9NWA9yciAUiBoSsn5Q0DVj4ZxUOmEqCHKp4TXBz4h4kOqmWRL6Tzf
GDm9Hq7mhlDqRbfJmMD1Nz0gcuTWiVPZWGot72ZNzY+RBMBg6rNP0EcaGiHepqPS
MzoU6TDdf6D0d+XYHpwZi153JZz0HZpk7P5S3D4PthLkibN+2z61PLdYgkrfpFrW
iy3/PbS5QHmopYiu338tAA==
`protect END_PROTECTED
