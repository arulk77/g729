`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+VXPJdb+MMQPvRA8NLgk6oayzz7FjN3W6fZvL04B9k+
/P/ZmgoXYAlkARB+chx0GdYeCbL2J9w8/XOgy9seR3OQ+nBgyAgzP6k5OJukZndF
A0AbnzABRTZ3vxhAx+GMKn6Ax5bGNPEpjuLYlNhPwaucYtOgUaTWgsP1aHXMTzE0
5Su+ch8K19Pp3TKAp8n6m26ewtycxEfcIc4bacMngcLaw47bjk+f842ozQDdQ5fE
/spnMBZBl5mZVrTgc0mm8x4XIxcYZfJmthpmNzp4g8M=
`protect END_PROTECTED
