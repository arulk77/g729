`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEDP+F2GLEmsd2lsE0i6SWsgIdOtfvgWxhoZuA0wPcz3
dRwisvaPxFoP5A9rl/a+Knjbkid+bH9HhBMWMD0avGKopBsANfb3j8or20YPL+Ru
OEyhnc4BPCrjDMqCEPi87XCT0BM5PrPZ+XPJxpSQ8yUlBqhkeSNV/p66nXv13tcb
`protect END_PROTECTED
