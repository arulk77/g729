`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCDb4AOTFGRFimlios/FxCVuzUVvWWTdVBVx7kuiSVTU
J9H0yzcNiSyi+7nlmk9EOkQF3JjtcXiPvBIeBitITkZ0BQ7xdS4xd6JC+XpqjcDX
zsFELb9sbZCoOuf7wRUc8SpwU0SdIFMDXO5hHf1sszA5Gz+Nt6HKKtWrhLXC1KP/
1RdykcVXN3281xp2OmA3dqIpkmnoG7XvLBLznFUCKwrWLbau6JEhIK8UoaWKDJDZ
MQuUnTAiFK8OgAmHt4B+z7yNu/UzTRD0itpPGxpVJYAWBjYSaTmfmN5jUwCmcZjt
Wz4Bkp93nv1M5H6pGRlnYJ/zYfJrchOPTr1oeui3rOv6CIxmZY4n+IbePdxcUZoF
`protect END_PROTECTED
