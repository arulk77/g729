`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBN6++LKr1sEeDFmA2MImAzlI1bBGkr+ni5Z1XUN7J/V
guK419xyMBLqdf4I+3x3ti8S2OwMqCQL2JM8wcKal6jJCrtnfDF+xTEdIHj8y6jp
uDlEaTebfHK1O3tACIGTrqKyFMmk9RAlfHnN5EAWy8KReNC4uGIQ9YvAsEaPTvTb
`protect END_PROTECTED
