`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/QS/yJ6IsIgRabxCW5ETZEOfn8QNzEo8/skSiIvNtIxA
5cF/Lsm8PtlvgSBHCLTWWHEbNtJvjIrISC2Xt6qMFafLtzqiVYyHbws6nd5IE2Q/
Btwvzg2eQ1RROAdr3o52k0IFy5d00aQxKqWSH6uHky+KDbc5Frn2VS1PqB/LH0OB
/ZS2MjkaV2W5ue+Sd36HIu7jJx04RIuAqK7QO0DMSq1cKPXU/M+OZEysUt5rysnY
96Iu5knsBiA6qreg2PWj2m9duhIFp/RjTjlbPgjauzApLg19ssdCexU4fdiT8LxV
cENnUD3C3uUCX0TwAn8i8C8pg7jsPIuDYG20Epl7cBRmJXEeX1xCDqIUpvX0aRj0
`protect END_PROTECTED
