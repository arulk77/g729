`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aUAz07QmwRdDhdxP8CoimeyI5K6q8202KZe1ixrfqClZ
hrDlfomV629cpAnfk9f14kVuMsREQ6KEbCifUKAwZXYo3Y3jhPp4g81Dfsk3gB9j
NDKbc2aYTqDHKOMVTsqsL8PaQk/0pGF3660s3rGFM7wN1o9Ba67b3LxbNk0Eubws
IRoK97UNZO8VCsTwtow6wfZzA5a4RUoDF5ZLbu6bMz+8aOEz9l+YKoVT/YWeZ9qp
7uiIy8Nm8TLgHS4K8hexlZUnUTy+wAsnJaJI3A4YYk3kzWwX0e5VCbx9Wfh/HswB
GkwFKDTN+i4Y8SUVrfPcXnQJi5fZpboJWfvhvKUrbFRfjlM6wPsod5zCurxVV+6R
va6t2ar2WbYwd7vdVyz8zrbSN5kBqahXCb8Xb+FYaNt+TWq24EmCvHyhqvaRUwl7
f9u5XyXDJCf+Jdeqm+HEirkPIF0yLyQwSji1vOsbEYgBE/Qb0UKXrOf2Ic16h1Sq
1IrgDsSEuHOSN4oAje07v8hOHyOTVValXsFrb4/5oSQ98XF9nKyDjtG7M43QRywy
T8TMnm6NcWRGVLTlTza9JVzeE+D8e8vTagvl6K6Ld1CWQ09KI/uygPMlUW6Xt12R
oj0Nobv3/UqGTZtTS3invwepiRitiNX6Rk99RHSCBgc5Izc6P3hyVxD1t7cdZ1dq
Tbtz5+qcN/3YUEYxTkgS2wxHMW1myWmNw43D6sL5oi7akqom/O4uzkF9B17fFcEW
rAaPPo1Ud/xfboHeUgG+Ui8dV2sGgNcxLzfjIMKj/r2N9gdeHnBa2LOIlvF/QLrE
SWZvJw9/mflA9r/8r1IInMZP4wt5PK7sGPoZrCJquQ0AMgcTpnsmOmC9wt6O11hv
vPr2NUqs0XaoKwF016A6we4evmmBmzSJ/lTlTikWZUdCz9hCdP4r5HKgIuZv0Tm5
D2AH0zNpSMeKFLR6kGwmxjpiux+XqnUWuOIgnAazLqX67xl3nsugmXRZafKheDWr
Lpt1LVKkfLR9irnWIOec9D2VFU6gLQTA+vpzQeZfx864VB66p0I6mgT8CkTlF+2W
vuzRkNMbexL+vJut1KLDtCJpC5mjE2v/EoHaAK2laIZdlPx/nKW/8vnUnV6+bYFD
42WXddJdEww0RB0lpYuzB0CYhISclgTs+NRPSTmuCj7zwRNFL4NMmYhp7ujTyqC5
9irEwLLxMvdG6ZxO4uFPmH1FuxrGkIbcnbGeXl6GqKukhIwkhYzrLvGed0SH8pZw
ATgmAcbYtxfLap+qDKElxITpjOehaclTQs/HkkRIhJn7lP95x6ZhfvYKB/BzzO9q
VC+5J+uHI44mC5ov2rBzglk/ZVet+ZxxwKS+gW592GzVNMIZ6hRhFPDtPWD0b/Yh
Ihs8oWpfPnmyES93pkY4kWpi12i8VxoitD04AhYgUO+bBGSGLM5fZ7toGHxOHgb0
WRNhemxES1zjtygNLG5Ox9TXs3yQL5kG2oPFDaQBxt7J5jux+nCKwN8f9ZtAcU9h
ht/JK9T5aE+az6Kj3/z1qI1oOxMTm2+F8zE9gvh+vxByMIDnZzkaRVMiXvHry69p
JwssPaPsaNoyTOwNFJnowXD132BRWRInReC7E78FCcjRXgw+6lqL3+/iq5XgvPuR
ah3UE1cZoTSSYII5yjJrlSTKBbgiQWurC/DfezLt0oKRl1jVXtZz8x5jv05dr/KX
UHTSlwXLP6bhKv13qkHuxob/1yjGJ0tFiVTsO4rFYF6q8kwq529ckSAtD2vDMfJg
ZU38PxtXtCwwbrA/tUS23dr+Mh/DK158N864xOoEco/KrYfF7AzfIeBFMDVpdWSi
36HtHJzT4lHJl4U6DW52EB7o00CEC0oRMn1nIyu16Deygsn6j+c9qfDu7Vq73bLF
R33ws9xW8XL3f8CnSKqTcsl3ppgxLTxoX9LYWaVzXmY4dQgxiGm0GsaI8yjhTBhl
JIpSseosH/YNpHZXzc3Agj241otTU46ybj8V4av0BbXwQaOKzr20ACOEa6X5zqPD
Q/iulMC04kGtiBbTdilVVOocrpjcNf4QASOL08o4g4kS5H4RmNX7HHZqsSyUpKni
at0bj4rlAXTtfZ5ZpwWyY7nb49noi+NXsxGLkEf5OJDVuufjMTV+0c4Yh92JbOrF
2l8zt1SIV5ztf902TJSlBWXIE98bvKyNxwiJqluFt1X+X422o+6+oYWQ/Vv90YbO
28WHAAuEH7b2lykO1fCBnOc0a1mjPYOEmYQn6JhcxaNgwH3UsykuoB7hicYxtc/M
IYcgwp+2BEqde/P/xNdAUBG7P0ON1Tql7GhBEZDdMHf4nkP/vAT1JQJzxvnkEpdx
89WiPf6GnjGTUSfSQTFXKY8OV2F/l+j6E69+r0Bdxx5UhcKAYHrN4oCi1+xIKpVE
awiIApnF0LoASYKg9R4Np910btvo3r7soi7a1HOtE6h6s3HS4odo2DRQ9/y4r/Vv
sa+YdkILu0IfY/KKWxyy0ZvGEyLu6y6reB4lVqvRQioUvA2fWgEEo6GSA4VRn5BP
tZIsuoD7bXQDBAPIoz/nOqxHnofW7yUuujWfcOt3xyOnsBqwm4+OPBWQ8L73LZ5h
CJ1eKHB4+1NXehPsV1iPzalsE43pO9FSuyo4bdq1JUOAxXpYL5qd4GJnHe1MWGyG
kxMSn0qEw9dVD/EzoYCdotI0YcZD10wQHh15y57WF5LxBsoV8bYQTEAnjliRVIxP
q1EJ2HSjciVHYsc/w0V7PG7hd/SaPuIu+copgk9g2Qw9mD5Rz4ugr02oy5tZGBIE
1l56XbW8Z0F1VdMq3eej2QkjdRo1cL4+MWhNSz/0dvij3N69jPklMXfrzQJw3qUB
xEi9IAEW2ZYzW85ceLSmB7p200UUiDyGAUHHIZbXus62cQIsgQKOplb7q/XwmAgg
5tyzvFrN650XHC4NoNsaNW8PghmvaupxLuijV9qBhdBo+vrStp7J82M6ZlDBu9rv
aqO01gCJBlJSFZBDq1UIFaM/cXlsx1aIw7o/OUOQQkLTnwC6yNQxAJBPzT9RmzIF
9Uke+3iVNz2k6SMA11+3hvreyNpwWA3bR4upV30nbte/pYTOmdy4H+q1g/7Pabwq
PVKqzlX3HRkLAx0yvdfYn9z2IMuIl2R9fwwv8ipxUGjHbqNOPkHmDdjdmY+yflxD
OiLrsE4b0u3iibedtib3yjFG/edpDHpIWEwsrPDE6iL+xAkkOi05ze0UBNmKa0oS
/kds3NuJyy0wp/83Dwlgouq66qFibt7CqWoxmFbaPg0mNQT9NzUyRZBP3hXQm8x2
q5h7Z4E1Cgg0A8n8KFqWbormq3/qaoBeIuwoH5Pd4ljZ1tAul/rSXsAdc8V3RrbY
GanE+N2JwumrVZKlrdLUq6uw2aG+0imaoThX7SEcV5y4KVwTm/C8LbHkfbmGsGqr
k74wKm0wfVPfS5DiJ7BErO1S1VACAOFiYSkTFulgV5Regww6UsO7sAIajHhR1EBy
A/RUhQYXTChm6HRUMhin4K3I3ttvnlobTztsGnLQ1G2n8FXT47XLquohVb84R3eh
Rd9iv6ansU+IjpMautlwg7UeMgX0PVcqIGsy9r39YGPAJXMLxOaUq52j+eMpiRXD
Ee/ig8C0wckZ5c3zObXKxnZdYORnyp+VUK/2B3yZ18f995LRu2fzE0kaF5HKhlIy
ZgMPkEKB9Zjw6rEN1PQyA6mDkHfb4Y0lNDiHGzJMja4hoZt9OLySmqZl5y3rkafA
WiwqxXgp3/UIoaKj8sDupuaIjtcHYkF8GSnpLcObj8Nevy9WjOV9pOX73ivtIV2U
5EhLzdmfcb/lzod6q8LKvjIKJ7Nc1GqiMIktBVtHLmH687NPDMyWbx44jCL+SI3Y
DCaI/nEOk4TpBBgmX75jKibC2sDwGsvb1rnxRNyd8+nQRtNnpTnKmqjdifdxuW7+
E4aOduGAtVhDI5eVno4Ah9N73UVo73W6Cyhuj5s33d7dwtot2GmerxoU+HKHNZBC
ysIezihFabKfw6ibMUnca0Tw+fXmTqV/CS9zljSPCRLkBobr9zlRnvwgoLN4jLKM
pMI12Jw6kC99vISqAv+VA9aQqIMlv0RxzVq6P4vYBf7W2a5YxFdD83YAj6Rjsqkb
cG/lwhJ4BnKdiJNQVNdNP+NPkDAUeerKqCuwB96ycpsLQiiUZK9l+NKjWl84R1xb
yHJzU5KG5ibwT+ysd3X4wABkH+j5eQGdeROj9Hagzk+jEQSZJUOdjVGyr/J8Eo2Z
u2BQt7JjhqssozjpydGg7LA60nEAUaigOKW767mqw37javbAe8pSWftBx97KiSuT
XN68tc9rcN9V2aCpBOzJjHP7mOhBDaReznELhMjcVSs10hpjtWX3aN0Z9bTJ4pFc
ohok2fLcJh2587V1HVfi7vhw4iWsxXNJRevBn5h/VJD6qRrsBErsDQPBgqksz2AE
MDNDLV5nFSWKjrfxs6+h+sEoE+YE/5bmycK6+bwI8xQnsck6qpYDumh3fsG45kgV
a7LYFH5rIOEa0T0vFN/Jlkrm9bD1OOiDY30iq7vLnOmY9grFkzMXN5roHyBVAqG2
w36AUW37IOf/V6RoMMMrj91UmjLjut02vT5E6BQRHour6VKIofJtPtUY1jM7avSn
xEnngvRWpHsFqP/7hk6qhquMJeKWiVz3y5dI6jfqOtmSgXNEgCodsfqgzMQsGDQX
QHsr7tyq3AM6rFRCtdB0KqTvFKBWyJf7nTeSH3lnYQ1zLdU8fe4sCtoV4NKYvODY
apEnq7iZonzHXHj1g7Y1gmFXV92maGe3ysmmdMreq3o7yRfUjtots2c1LP4Qo6X5
lIQA+G9nclA2bjlBTNIXi8PIHOM7/U936r1Ei4GStYHiuILEm8wmBAO5xZorCODa
RjBM/JaKgCAdcSdxFEWmIhf+fPpxymCVZqkpy5D43Yyu26ugcZrVtPgPYGpbZF5S
Fu2JKHag6FYoCE0upepjaMdjvLJDd6PehUo2VEdLvWpU73BELE84TsuTv0cHQmuB
FhjxaxMjN+tG9XDk+fv3B7cM7WECcQuwXHJjUb+/Pp9kSyjP3ZmVSKkZdk2WELJp
kpS9r1Zi3KVYQIvKnjByYaRiLtqvKjYB1bg6Hta9Xd3wUZsYEMVuf/rJYYxBiG1m
QDXtfHVMiExSRoRF8WR1gJvxH0M7ydPNteLUHeLkLzHbNqyuK6BiatNuDvscO05W
STfmuijo/oGRkdOdSZHoWTZA3te+f1cKEFJGUVw5Zb7UpYpfg6xFGpm1Y+pvndIR
Yv2OghcwCCBJRGW0ggI9a2YVK4rGcSvMp7q7xm+qh/sltQYgqEhaAFANK5KmRmHC
p3rnlJjzBdt4Vx00bc1jq2RvePbNa/vxZQF0ztAMIO18nchGSuwFthTxjWUMVxb8
ghWRlti2yKbnyLl+4nrYpYqH7BiLvGR2eIj18LmDrpBl0cf3BDj1/oqv4nWcDPYE
V1zvENRUFBCrcYA2gjH92OQDk2XjQLBrkLswIJj/izQmTGtMKmCc+DMIeg2gkdef
hABxoauBHzmjETz9bd5x2UlMZzdwgJxeKx1luZP79TzTEEx4FLC5JQbdqSYzJeH1
gPzcdfnse9IEhxqc7CX9c0FQFVDWMPh9S2SzoPYBchPSaurdhl/kYlW8LQjwl2iS
HuJDl3fvTy07vkF9D9Apa6TF6Ygf9HFWO9urXKwSVjkkVW1JU9cjzEoKouU12Iik
H8OJGxWtobN0lenBfvMySivcstc+VyuYnTk+PN59R0BAQK0cX/rpqPtw0Gzd/Edh
s/9p6r43AfAvToPrya9/yJkyiwzcAKDNKFeEDR+mJ3uGthagebBAWg0BbNh2Hdm5
IgPHyLjx0mBCWU4/XA5E4NDQ95ihoBxgBvr0Emypo9KUDkFbZqaaM6z6o1aq3b7k
vUagdZwUpYf9lXiSjpHCNvMDsjhn2Yz/LMdA3xCTyM7Ye2dw8sSWNyVO6YM+74j2
nFlIbVGrGI6b/czVJlVLpJoktpJrww6FVQaGsVbMenBoJJeYYSm2qSUsR0HjMqsF
B6GGKSmQZcfdjrb/VXHq99CnUk4CnXYSr4xY2SUkoCK4ezhM9fTpSLHcWDv46K8P
h6sE0BqXcsF5pStmipOhkVxczZYkfEmBRnfkiwnZOX0B29eUlifBBwnlEXOjxhvQ
f4oM/TCMhBq/dquXYRDWmK9Z1S99YTZUOZsEBjeAaxwEuz7h12VMU9XhJXAep9Yr
vlAh1hPO8rUsqhBpcrBrj7VKMEoMk+HJkqRA++Ai5jaiiNMISPyANeAouGGvfIIM
FupyyXgKF4/ICzpFn1WrKJ5xKgYJCYivVbm6h2lEvykI902seoyJjJ9zZAbTRJkB
lZ+OmccfvBXBUuQdY+h60vgYfwV2U/6lcqTtwHGFD66zGv3cu9P3lahiR971rRcC
w38/nHyzfOJS4fIDECx8W41AcxNiDuWms8jWgeEDTfOoM+YSP7JN1A5FmaFHGF9P
wy7e1+jOulDKBpt1se7iO/qTQr7NocGDCq4+Exc1AEFPkvFmeu+yFdkHzq9ksxfr
Rk5wCfKx04fUM4O/2Zxr+OPPHBYg5yNBUHDsy1vuvPTFY4wCXloJNQP2g4jfYQLg
5z1cWD/gP1stfyjCDc8mlLyNy0tQwyk9zmfTXUU8aVU8GOdWwN/1O1JFIu7I2uE6
Ji7GiCZb/JkzkwWg1S0VTtuvRVlD2dWLJzIpK17J1PDIN+Kb+6h4rwN7lPgKoJ8J
qp5qJZS7uwBAg+2gA5tx/aqRJc5DTLw43oFbmyt53dTp9+ZMO4Ay5EbslHKbyHV2
geu40/DlQEFi5JAXlXydy6crRDLUV1vwf4xThB8aqQpRtBwstmdHumhXLHXnSiOw
dB5wbBR57TYUBwyjNTpUiAseDYPqtp+xEze3bm75dlIy9MZ4Y6Xq2bHRy1QIc+dv
9WcuaCnfEQo8o7zrWmzEseDsdogTjV1XNE73iS8o/eFsmKFzcWpvBU74yhTaggmg
ey4e9/HmL61ytKgTFYIbBkGh6j+sGE31esk3W8YEYtvwiiPKoJ7OcCNv0fE2tVo5
uj9U4xLMRZt8Ouv1CIZxAJW1f0B5G35G+wZM6viCPTO7FoXuLi7Ru+ZXfj/Cxa37
W3Bioywisp5NIAAl8MxqimtE24aAqr+zw5viDPXNEcKIIOhBchS81QOziMpiSEYx
bb4A2C8/o5yitIMdAjufPcRaQTy3WK0xdPngn+5PgXKxjV8o34iikbE0otSqhgvS
QzZAi+QabvtfBagmeNGEO+7sDAiQocxWi2zYLNsXwEzRqRgArbR3AV2/p/TZg//e
gD+35jQ/xp+EZF2lWLdT7Nj5AHFX8MRZRbJMz50C5UOEQtx4jJhZGGW/WttaQr00
yrwe778bHfP5DOU5lK4JMXc6YauSmUDV02QRPq0dVEoo2zvlhgNPG1B216Am5LBJ
U05g9XGtu8N5q0Slhs6/UXun+9croZOxe+0mWc1+1mIUjhocdqnjpT/1vl6ccsbg
/1VPkwyeyA16JoZZHi41LxBr6rqku6Hm0ZJkTCR9jtTjfCJm3SvxXRkcvoDXdDEn
6cHmdVmQRts0vq3D22v20DtQVqs2AwZ99E3eHdPOSE9XZM6lQYJQ+hegOJj/Gaah
aKcHTLuAytbdbJLUSctiqdobAsiLlcQ9FnMAv2EsZwNcCHp8e5lDm/sJyD9vSkGy
5jYqklMqGwWA773mGwe+k/kFZC2PjJ+kS6FJzdZBkba5Y4RhbrrDP+i9TgnB6Puq
FYQqs8EtBaI2aYB5E7d6dWW9xreBvYADnkk4GYruIYAscQAohPHCRPQneSsmg3UT
9Q/6UNRsM7AMKNK/CTBG7ziqhQdL/HE1bmDPNlRNGZ3qnlw0qvHgKGq70zld0hR9
8X95xQiPzCPxsUWmyH78nwXjcLEly+eUvkZpLcrmoWfrbTId+3xpUZp9K/Kk2p2u
JuwB0S3LUmGK3tBrqHjJ3wjlPl21bTNfBtcRe9+rXNEp0mXI5hxuxRexyFZXjebM
MiJ+6woJnzPpFD/1EAARDm+TTzjkHQ8KiuOzxpCGUnAgxuVCDz+YJigj1z1+89vh
TW55QMeqmqBtPrGPGW++542G6RAWau+YhfOJ209qm+Rx1NQdp2D60CPnJHx+dVrc
LLjtu78MN1M2is6snKlBV9vuWUjlH97A0F6DINKgKyDpRPNTGwIU7Krf4y97w37o
69nd3OfHaiEteGA8uDFCVT1PIBcjmvhsJmOfPoNAXiPOfv4eYWbacrOFZSGUNKTG
ntXoZB1jf5JP91vOMptdYTrYyIp8Jg4dul6l8NFM7kjkdKpWyO8ajFRTp6sG3L8S
8WcAXL3MRwa7j+EIMayzzDMBNK1pwpD242iHTzge5a0pV+UAsPsdwltnLCgBV8Vx
9N2T7rvDe9p2d+aMjUeuiRHy/Z84rqkj6ThYRJ2LijRlO2VF+CxQZ26/DeougGf3
`protect END_PROTECTED
