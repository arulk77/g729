`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CwRR5v+oOZGErXwjR1oTXRejf5iM2nM+uaP8bjEbPPow
99qeIH5sPU1R5JWy5lpYL9JeQZlqPJEKg2AakxANS7daJR0TO6LJdi1ZM/XZAQrA
fM/kFFdDiRoGRhnvDdXnHE3WMQejf89BOm8Xr+uW9+mGmfuERDAcTVOZiKc+CdCW
pe4AyFdl6YYv8QsRW8dRf7HZBJzM6WHQJK6qYvRYTDr8lJJE4DEnKUCeOBUFxNjC
f7LNIsJlsZDRAjeXXlMdYwlVMIask1n9fTgZDqWtqSA=
`protect END_PROTECTED
