`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDqyvtQGSpmHDv8zTh/H6ephMWLEn+XVpTagOguaGawSSc
9jVbN8E6dDO0wGKvZcFkoJAF93M3lI/LjCkCybs6bzOJfbeDjik/rNz9vqCQFiJR
hi2ne4MZtBtCHOK2TKS4+mkcBjkSMs266AXFEss97v5Ce5SaNhN/kkSvO+/X5Euo
oLfRZn1p0YpwByiKIgwhLqdKcCtCztIoiXFtK07cPA1+R56Sx0NibciyJ8lRuZne
qClLoNvNgW6ZciJhLvtxaUdO28YW7uCfWBQFdU1elR/gT0mX8K5BnRcPbtuhyjN6
`protect END_PROTECTED
