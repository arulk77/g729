`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLIj7hyF7RSeKkIQXmptiOxoX5DkZjpvsa2FDI51w36j
2rqDEmUEOhmVpmS3CW57Ns8ByTI8s2ket/1gcGe02esLsxI6fYu0fKvVBypkEOTV
KhUaaJZzrVXICDaBnQ40YZ2MZGMwRlkt7Ij8VZuMdCBWL6NQOtBmZ3IheTN6ZHkC
mvlAP8eu5vmDhTwiuXWFU1YUJA1HEfIOPIT7i41lUtxS6t6WIB7c187DtsAPc55P
EoCnHSKCfk7/VtUxexLc98iJbpVRY5YonxoFSed+E56FKeosl84JDI5JxU16mk66
DQCjzbHgBroHC1dmkn75SwB1jUa9avNkLFVGDDsrcLuO20XxLPW+IwzTJFnTmGvN
`protect END_PROTECTED
