`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47oWCwAyJyI9dvssZIjj1N9zB+ecJqsWDKrA0lxyMSZF
AMLU4bEFHqyx74yE4E76UUZd2t7d5b8fklPPdBxjtiof6AYnGAsR2p5wAkWRSE5f
mtA5m3VieFGiokHSvv6hqWCctn7jj1934egJIEtLhdWlqoybHaCWZMDsIJdpHWXM
LU7SqKZhBxxW6bD8OhurFlqk16lZ6f2K+2PQgim5yFO/0Q0PzJWy8/WvnVF49Voz
SfST/Zt9rz8IZjVo8Q72MrTc2W70ZsmC2BgC0NI7o38=
`protect END_PROTECTED
