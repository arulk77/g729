`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LyBF6XCTpU1GmFmj5q9bGv7jCiFl+RsBCoTVXV2+wmSmbsxrOA7Qy7xBTeFQmsLY
kQAYALTL2LLNKUkD5AQKcUDTcLTGM8Se8U/PAPZ503P34Vfe8LulFu6ixscfw4u7
UeiDTODHcW/0oBCG2+DMkCkT53kfhebelz94w8P8j1AP6LxeMpVHx9n2he3PP8hM
YDB6P5mtycWn3qVqhmojea5LK6GjwqmI3cZ8m26gRxklaII0l1kf/PI64vuS5Yp5
mSoez4KuxCXReORiDJpoLju4d97p5hOPvW5dnTaT1kwDwOiFksVfMghldCqKNjaS
M9ZeR6izxuIETPITyNNn/cQygMpMVS9rJYtSI/B9YJQ=
`protect END_PROTECTED
