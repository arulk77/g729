`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JhFUYKU/WPihO8G7xTFUQjL7FtoYtpWjzYOMEZWtG616ce7sQsoAFvBZFofD7cUw
S9uf0Y3Xu7LsV9PBvjo4jEOKLqCJB4CXJxY18JwrEH3JP86bAHjf0JyoHk8rlQlC
ki4nR3EhX2SdiUhPl1gsPJhMyyAzMfzPgWFLtTyHm35Q6hofkfaYjqGhWZ2y5feK
XDFPCdC0l/A4gDERhhzCw+LX+DUT+OSxWgRUe05hDD7J1b8hqv/PE2p3VE2WFMDM
ANNBXbzJoHxYGlVXQTKCryY1BfPmKJhYaY4vgeRabge2/RFjb1NNnUz75XFYgzS1
`protect END_PROTECTED
