`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDQgTPqG3/CllBZ5UJVccaH+WPqEvET5ggsaUmKe/AZb
Do9o3dK0bwinGwJWrebNiE5aZy9YLtrf3hWaHj9WHt/hESReFuRG3AH+Lda3i4Hz
iJONpjAKVDOydKxx7M3QsTA3rrmMPa6DuXkgQ/HzF8KcSTjnxWVI66+4pCYsW0Ly
jKR/0exo/IwugTMjey3En2TSfSpfqnqz00Xj5M0cdIXH1CdEymYf+35ie2eOlSuF
xK8HZxxnM/JZuIBtkdAHgSHxBx/+E6jwxdHgE0g85RIo4HtB7TGGFb31eADFZok3
8//7aPmVEEIv3Cpg6Qonm2fsKd++eTva9AsKRyZfKQBP0JkPXRRYSvxlfY23Pswi
BhwCzB2cFvCAFg/AAjVNci9No1aKQaworbWySfLkD7+qDcfVZ7Uh7qiut023kSxH
yA4U5gxp8BIcffxyB1V2yQHbYjdeBdm9/lUptbucvAAQzQPfJ6qaTBwZ8rgSPSkd
p+anW7lbQAKIsuPvzijBR9gRBG9e2Sv/bCF/Q3ykceIco0GfsHIpC4NrhiiX4Zax
`protect END_PROTECTED
