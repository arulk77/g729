`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIbto73aL5faVwH7sZw6lb23HuHxwfJnHfPgsTh9qX4g
/n+wZeELEKnyeGmv4ry20JB84El/wOFUIFykEA+mxqGd1SjFMP5+URRO5Oj1IIPp
sY9oiS+jyi4oj936tBhLRUpPcprHNqREm6cg/54FfPBimsxGEn3UzmE3jKj6eIF3
RbVZpbRzq7hXEf5tVHDh7qXacZ5nKufQHHgNlhzPkhM3BRbs1uk4pzU+bfLkz0jL
rdW6tlVj2jnsmIl6BaSbGrndYsjWG+EOn89Sb81JtcmlY3HpU7njTduqKimW4oEL
jPik1u7vJPH3i3RIedox43oLI+vJ5gbxPOCr5ksC11l5Lqs6BLWuTUl56HAyFPE4
6XVnvzkNZ2kxx9LkUMWxUDLXxq2QqQ7hdUVE65PNIUMGraaHQTPIAEZrjghcccjV
US2x3xtBxEcMrunm72VsXP/mtepXhF6Ruk6PK0jF1SIxeu2T5PR056nzjcXz2pO3
8g/9PSAVmKHzDWihKonYqB7t8nAuA24zt36707DwHfhra6OLhhiLg2qtUbT62Wgw
qiN/p5PeEP6yb7oU7Qk10QXwhXMyvcOBLH2qwlv/ko/saU+Vd+Z2f47U33ItLOTZ
`protect END_PROTECTED
