`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44Yok38WGT0wqLXYAfwXBAUrkWd49bZKWaojURnyzQp3
Mk8KpeadkWKsUG9UXVpteN6PSkKcXV1gL1d01jJQq1/Ss2ZxQ0M5pXefrEV9GuLF
pnNqpgMhRPjyyvrPDu2bQWBUl62LT4vosKlx4cPaxM7eVB4p4E1G65QT+dVYqauB
bzpXu8qa+YpOzE9utCzpn62sCuLGenhHnecshvJhLULesGCxKVcG5AmxPR9xbcg2
96YNBODqkRCNe+i4H2BbyVh3CkJ5KIDy3v1O2Rktaf0=
`protect END_PROTECTED
