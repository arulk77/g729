`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+3hYJPiTR+Mx0jQY1vnpr8Vk8C4DW9HP0Wcq/kq1M1CTHXyFYzcifT102hbEdYH2
8wpqJIlBkRZlXJJhhO/pX4EMOuYhsnZmIPRQRrPsn1lCUwNQTvts+j1UssAmij5T
ebRLNQ5FKiT0vTOB4PgLCIreCB9pri3E/7EHRrAw0YSeX7d7c2N39ejbQAPUcvHG
AUNni+/0nUEONJWzjhrOTAtQ0gyG2izXGW9y4qQrTqpv4wYz8Z3gGLXGAQdx8PBf
ggzsrLwaZHAW5qM6fBn1CU8Ic5BCIfjO5zqa8xy6ApU2ijBau/3TSvKhKvLCafPy
YwEnlrvUT0nigGLKAIinJeeBe7nzI7Z3gUIlJiK42GIh0wRS5ucj0NgavuJEoPxN
udL7JANP/U7OrreUZ8BPZMUa3TxX8bAvdjPxHvOHka3Q6cT/YnqZnIxJOQJhwRlW
GLtuWVvo5aGfZN9aEoM4fTu1GdHQzz7EWjvVo15gvH3jjAfnQCGDe/THW+k7E71q
5mDL0ESJ3pKfn8VgoHlxyGJwO0m5UM78zcE3AJC3ZKD1PC0HnzIrIPRNkMi220r9
FbRYzjgcSnZrYI6jLNPHcX+TEivLJ1UvVGLjvFZz+ndt9mstKf3PLz0cAmmCLnnL
ppOLmY1royk0WJtyf60Ag+NHvRYvK3DXQ7RW6akYHSJvQUv9TYFjQqqor2//9+zZ
U63WgbTwzH9TTpQzupiQ7w2w+AcGOfz9h858XXtvC6wqS4BW9GJHLl/9rgfYh5ih
FjUWphgzqxlKHjqQ9lN2AfMSBMuA8nUMm/G3D2ptkXmNLLvhmmAONfdrc5joN58/
sF5OM4fnVZ4IJNS+Uvw1/xWyXSSswpMUInF8pR3j2QybdSSrNI8Dfc43IyZm9El+
vk9CRp/CuDO/8Kg8XgaFmGzvUo7D56O2c7jtJ7yL09OqpGiwFx1LQCNOreMbMtJS
Rrv6hkgpP300FUZBZncgnIlHSWPB8A5hs5L+nZSuo9Hc/univZQbrNTF6Am/w9xM
6maMIYb7cTtMEXqnkJy5dOkvDzGRf6z6grW2ARlW/iwq98/YIUhKUlcmkMI0GFZf
Yl2SGEbhA43kr0RgiazVu21vmcKHBUVxPKMKSu4UboBp9lTm3qvKrZvNnLBJt+wy
/pH8nTjlHAxJF0DmGvspJhZrMWowXT5xkMB5rcmnZGJUq5IbmiQPKcxzcuegBsJl
pxUN2Osz+f2hUnHQs06nlhtkYG2+cKm+0z6AuFNn1FF7hk4B8MazBcY3T9O76gcs
TM5hqPtiAGKilF9HOPDLFo3lYXrVzb5p14cEjMHy2iUTJSh16Sd5Iv5TalymAeRM
7/Es2aQb7OVGarEfgzpFHokp2be1RvXk/ezIMyojMrpYhBMnrJtAgzhaFUghlxLn
vXwzmueLhRBXnIJAcziYzzD0AlxqeHSJhouLUAaptj7Z3gxV4sRPiBbvUdPFtxhv
CA6729BG5LppGsUR5LYE3A+ArwAu8HFuBnZuRo/GzzJtSiyeIfqXb0CvJ+L4kfDr
vsfwjc1GllukRnwIPocwzzkDHyXxRAFb4ucxcYC6CWDMCoRQIr9Zxi0ciSvttorY
`protect END_PROTECTED
