`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL891EjRQDI5woej/08rn0BDKnx70rn6dWo37No2iwf1rE
uwCT4IDKQDe8P5EXOIRBHIpbN4B0aeXVS99ziE+/n35fbXsfbQvBB4GLpYeST1Rm
yUXawFaKiohJRh6cQvFTkK32QtatYMdmr2s63Urq06Fj6Fojl22WFohT2HZnzaoO
h9wXtqnd/2P2cg1jZxc9bPOL6boco5k54/+L8+Oi38ICWmZOy52fZNgNA/AjaXGu
/wdaQqWLNGOUO9E+jxuA0dT26D7tfJMCtaz2szC/6aLvKVUBbn4L74SdLnJODSZ5
MJZfykit9wlDMlz6lqUUZX3Q86gRni5qUK/vLjdZzvjyCniH3k2xSlE15faRTPc2
99W/hDyfdBBKIV0R81BX4NMflA7T+EAFiHqzOnoVGETtK6IUkQztf/ma+G5ylsZu
+seixo6FnWoTuesrDZ4Sr3t0nQPm8prNWt9PcWHvZVBH6MMwR9NfOAp6vHn92vGz
eyuZXNXyCkXmfX42SLTXKh0jLyR+nC7UQALgRE5DLfxlqj+z+pNQVO2MGFFx9FO6
+bzBbeLYRr0rbRpTG4SoeqLSb92N8WNXCl6IN0zTS53la+IAaM7HY6sk5VuAaM1C
uZLgtE7A9AGDNfk/EQpCiS7EoBVt82vMI5SuoM8Bav6v6pVdmW6+PeVtK9fIkq12
XGNGB5XOgmgDDGq8+RIwcLCqoDYwJH21BEdqlypJO8sY0rYeXGhLHW0ZlVqGsykj
5OK4Jc2m/PI2Q+jwCee6qtoTJuJQXFbF8Tw06WqErBhCqXl3rDfEsi21kRo8I/jl
o5LDZ3BLsTkNa/e+1OaOfQnW6ArUclpujbOh2gpvKQenLGTnefz38lPgdOtOLEPY
gpooqUeB4LQZEOlgTQqdOxvJ9XJHfoShfia6xQmghQ9RjBqfOzl36oRMIR6MYUMk
7qc0OGzoZ/tL3bmTgSXYWUm8XV+OEEYLoy2elbHTdSw3394/WhVqph4QJ2JW5IRi
vSR0UH7AkV5Dt8T0+hY9uY3JP6JJXt3oNDE1USL0HRz5AyySfavqQtG+dq9pLq7z
5JC2Iv7QliNZ4Pgqd5ZlRjrtjue4Y8x1zQVAWaqaQVVmq081dk1ujGTtVl2xOJUR
1HdmDiXUVhC4y8T2J15MkviDieIu5czTM7eFKfinOTZAx/CQh9RDp8WMbHeUhHaw
sX+Dz9Yro+dUrSAOpeWMjEJVFCnZdAPbsm04IoAhdREq26/lrIx+ReamWTTrNkHM
Z9kQzy6bhxxLTlMlY3LtwBcATICk3kSI3XRbmUCqGJJeSUUfxikSJLa8AZy2EH8M
NpOy0VZwsay4nwXxxps2Yp8wmh0c0KX6tMpN+cxZlbtVonGhq0VLzxrDHUuF31Ua
aAXhlzioUqWim4nDlm6QEFMS+VT8lIRwyP2E5YlUOygL/5AUKis0s0egNg9N0MYz
mU/XZgnD6hiQVLcQx43kzVzZpxVY94MphlPKltSIzFzrRo8vHmmn6MuQ79S43JFx
sdC9kGpM8+pWjB3zY7T8AjV47L5Hl2CTDigki8XED96DEiukvv1mjjKlfFHLuRfi
DcKvIhpWig6zUoj2SElwJGx485DHO6Ul57sgF5qJxVbYnrOdc0kk/qrzQDUxYpCe
M8ieoUWMqV/URrK2aoJVgVKBOuKG4tsaEmvyjzZNyB6jfUAvFI1skFGNjrIrI2Ii
p+juztVyrdxrw70yOdmAnDkySRq5S4pQEzmbpD+KQb9WHw9/hae97pQtMTt+h5Sr
u1et1zWY4x4K8KpNCBex7lCKfkx1oLSwv/M0RRRq2FmsrOIhmRWfLjKRMr7TOhzb
HmVx1VOLtH7iMNtwMgc4WZkPNC5ycq1g8fLF6C9/BxVEXPLPkPCvD3Zk3W7WYPU5
uJYPpfD9VMAjfQ/mOfYaGXXWtAMLdL1z2h+wjDAPf6kHhZq9Y5YYsi4VhAGfc5dX
8NxTvm+CCsphEMElY7jPC4b2owD9Lrvpn1uLRoiaUqE=
`protect END_PROTECTED
