`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46kA/+/OunimAhmHjrRWBghZ4VgizsiHoFVJpa3XunDr
UNEy5MapekWklmG+1niuydDWIKdZLxAEqGLa0AmXvNxMq1MxlIDjhUEKXZ0Q2qHq
Xltkav+3SBzluaX1DUpi67inz8DMgo1tVRiL/lUamfxVNs2Z8ksy047MTtfEKulC
pgsXjRphaeXdeWyzZh25pPVmOqtg1hQHCc9SdFehQ8lgbqPKHE0nuXslaGtq+YMg
DGD4qEwvKg99N/qfjYFxyh0cKlr3gmc3JJhQ4JdGvSeSOxFMyK3GuHOhjq4ZbEMr
ZFCTtlfTSNYReYmeeMzOkocprr7frQFC7rPrSt3gGy1+O5TIy8Pp/gB6nrHiBNTS
Xf68GaKxKaWPrsXQSUrERwG4QzAbi3qZ+EtAjf48YFpE6eOSdoVMh4Z+uxOzd9Ef
EdBCVhfvWO18k3PSWRkZtXqJHg3CYm9QsThdLXr46bwZuDNjPOfFSGFrWae3kvJa
nlV+yyQgHSeanYLUBsUvcmBxATKcH8Z4e+IO7v1JzgfiPxb3laE/sSD5+Y07jy9E
XiVbd5KDf1lEZM/5il+kTqtgifie53QOdyRiZHy4EWgAltZhp1xu4La3agcp8809
`protect END_PROTECTED
