`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49Z5O4IUoHcng6K2PUHO5yg8dxRM74nBFsCIvEmEmAoR
xqXgunh940HHxM0A7ETOlMej6qBs3yBHVTx2Tjjs2BhXWWl4bZB4J691/tH0sxWo
Po3mUsa/mkoF0xx87Mg7dc3dDqkIMYeTloLqBlskC3Sivkz9/+Hp4vdotyBpryZj
kKsE3jRRruQf6R+1ydUd/y/OhN+VErv2okSSHgWSv4o=
`protect END_PROTECTED
