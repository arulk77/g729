`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCStD8D9z1jBunBt8fbAmFJJ0qFHVu6ATR7qjv8XZJ2S
N8zn7PJxoPAGtOGYgcrgYsbQN3mB3XbHxPd5Y7RAC1Ot+mJK+mKBRX4y/u6ocjFV
94cm5y7lIgKvbcr60B/Dbsm2Dj66yd0pA6pcf2L0Rzj5+HKQa4xcwHBNu879JKGs
cXLR7MiAch8frmDxEoLxiKFw3dkH5QcszJvuGDi14WfXAK8hhn9psRFWKNs4KjFA
/i/atf6d+6aY+GrkD0dITizACYjH4qPKZT/CNdPt7lGePDcUcbZU64RrdxmFLlBc
xdASqeKGqUZlT7jr7GD3a9Kdk5lqlEm8y0yAYQFBRvcAPS38Xeh0le0J6Md1VtMu
JoIDgjMWHT/7K+pAOC4PpmGcOIvGOqR3bcJA5F0gxamTMj/9oqp3FbEzPEf/Y5FH
tCaMHQsjmYTAnWYr2m0Vx9cLQ5RxZmz4nkDOeGLuUZFl6q95GC+pOae3KqRbOj2p
s7QqVCABhEcSm5pSUlkFuCJ4KpAkjvDxYYB9D3LCNe7X9GCZHxXDLFitN5MOEhm0
e+njn2kxymhgqa5D8r6tJvZ3A2EMQWwIoNqiuOH4oAaETQ69T7VHpTIas+nnPJyK
p8kSa/ELkaRddeBUQixBaAN5ATFssJeiCzGOatzkaa2r0p5dqkJVbhe49xDvvEse
wD7HnvBH3FUEMYnfX4grWl+0/GKAn76A2IdxRgDWwxkwvUQNuZeyH1dhEcB5XTS9
++HJikmBQsP5uJkLph45CW3ApBKGxz7tFWbQMV2MoBGTtd3iATP2QoncMYjjiyxA
y5UPDSgkLY+Y7p89mVPowPUXYQ5UkXaMJwMNYpWJDP/VZMI1rwTTem7a4XdA7NSz
D0aeZMKJLBQxqP4g1ZW9hxnD4ZZB2l0JZhxrRY/wSdol6qWX6T0PRGxfvj5fC7XB
jFZz+/2sNRShzrB9UpBKAF/u9/CWdkLKENwvAApXSohmtXMBPyicfNvzCgPB5NU8
kWZmpaxzm6x9iPBLzbOJmXndNieIlV9NAYZMgSh6nsl03ctUew+eL5EB4jEAeaso
f/P4ZnRVVC+mQKgWBMt8bfG4fLY18F2Hn5RVMfZ9edI1c1woNFSS71ypV2UpWpb5
od8Z+779Vk9V2IIk93Sn89keQhc2XowK0tJ4h2dotvt/ljrTsJNU5Q131chlRHxY
NA0xX+D1uelL29gggTO85ITm97UpNr4Rkv7f00JbgUw7hKQ4HkbGhjzBV0YWHvV1
nQFAEQ27T+qtbPUEb8OoJLlrjpoPIFmCQYwAtqWy9x7hb7dRVekdh9er8tDifxT4
B/vP0ZagKZzU0s6cccZzaUDEcmg8GLf0pxnz1kcDBzfvxnOwxag/2PQqzPphA/KU
WOqUyAVniv/wd6m4S4izCn5ZjISggvsUsxmsSk//OmwskDAOTw3N7crALwk/5IAI
OCR+whgYv3crMNUSr7qDVVr9x1S9gxYeIfD6j0nM+OkGZkpf0IhgV9VZZiqYV8de
X66MJUB8YU3BiwIprh2Hm1NkNu6IRI1k2jKfNz4tpIXDCsmLXf2Z7pysPxmors4L
P6SI7uvte07fDii5KBG53sMksTkuAUqK/9FMyTPf7CfvacRrU0DVx9MM8zdc+FHW
9a+a744ZnvmuWlyXSt+Jiia4uxuEEwrIp6yXEsifEzU5lsXRI9pislelhXyca0da
24mo2uZ0qiT6bRqcBAcIa1vl7W1VqTHmj1hq32/1HNSLJQFtRpVEW6tOP3BfETY5
WoV4Tl2c6606tjZ11VjhG7ERCsWw1TZjvq6iHmAkukdY9GfmwlReg0dLvsDDzC7j
0DgcYPzJdwqUvQ2hL/9o2f2O+pwe18ipPNfoMWHwINRZPSUrD7/CZbC5ldVFs7BF
R8o8GxssmKHmfkSmaPTnEKQyv/yRVuqDXRxYAGyNQENfRoZ4FEAC4CF565DAIRlB
yhx1FY9cbcIUk0FNkP721ZOupU/HRYX2+ID3ah4vne9U/UevQgqlEMMSgr295FFJ
pvs7ivGxfn9EcWd1n37nHpLsGPENPi9n9QwOEH3DCIJ/HIxKIuwqnxuRi9XOllp3
3/I13Qhytal1sDwq5wWYI9W5b+YyVp6UJUFuBq36407TPrcQu4Cy4FwHFeb3WiAN
3Bl3v00YpoJFt1T0v9/5UQOZciJ35sHucCcV9eSdfZdiNfF3Rzsflfs5EoCNiNj6
CrDSJKE1CQgfM0OusEkmql1iEC8qEonvi4DId6S2YnxGPnlqdbNu/KP/5m0YjEDm
14NinyM04reHQ7Z03ttCUiYcmLlcmAVhJpwddcWDROJbSRfRmX8p9thbn3Ram9eg
jz2rOXsnCJmMEbM57DP7Afblk7M1WsYqQpSR3vIinzWEQbYDZs+pfaJvENhUP/P5
eWi7EpeJtYicoVmdEe9Hvs3I+DcHms/Ee7KdP19TJDLKtuuefgrA+iVRD/DOHNks
w0c/I8m0fFXyWuYmaonow8wDWno9iUlGu//qxSUOBMs=
`protect END_PROTECTED
