`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44IcJB6Q4noJs2sqdH8gMjItZXgKzU8OMk10ijeV8aSE
9jF6qB6RvuS+ZAPtIg6cFc2D+SNDeFO4bpfBTwsqh1wHKKoNCGxRxi9NLsrBirc9
ipjvVcoIRrqd2RKScA6ErR84rbSx7gfGT9XGcY6P/452QyB1J2qKYU2yFUAmfbw9
SE7JdsdKbyN8fqpnKm+S8op+8gtVlQVFxC39fR8ai8IQgPmIm/inpD2iV4wLTpki
oxHjto7fPBdszy+eNCn8/iOb7jApHQfySoiuV4rLuEg=
`protect END_PROTECTED
