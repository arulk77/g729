`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHGM6jc8U+Wq1R2lu0AGOzkcThDHiT+upAG42rk0oV//
rjReqQaa2lheSND24qu0EcupzVHka2mzXVKWI/2D/K4v9PXFm7SWM/BhA+PqZ1Fm
xBN+SSn0fAWaIGXDRyxe+L26mCTCAvqqy35B23rCOaL1YH8vTEYU8wErA2yfX00i
q1rENy20EJNcqkO9LXQPwnSKqfrk4kAcRsVggl9bijy2opdrrqQ+tFDDPqyI0f8B
Ro+8B8qa1VuZzUat5QUSalqUisntR8bqsXJsmEmMVKLQwdFaK7QeQgNGFV/frp42
Psj9BLxVSv38+00vljskDdcYmUO4k4OEuNLECUrYQjjyIgVllovb/4B4znS7LQHM
YT7f/mmwE8qw6GkvFV2eEpo/Fc8JMuPHEctjSwwx7Ec=
`protect END_PROTECTED
