`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
qMQJcbYbE3AUUCvfqngPYgWjzM249ASt+uQdi/9cnvz4w9HD/Wpj0P+dy3W0B9Qv
TEzwtgcbRrje6O3gREO2BP9oqmE4nIfkjKDMpBccwPqq47TVQBdUnkcGyzDYrxXn
ONl0eiMyKZ/alu98Zv6xLJN9WXeV9j35gv0oMC1OHi9RyNfEeH9XqVVzToX3ZewS
1zp5J+wZFMsRvKcN0FtmMVXDU0DYhMXCkBfMgak6OTzKZwCwf7UE4PJXnsDtP69E
JQoHZsUDmkQK/gjrNB8L1b/iPzASh/HX3f5HJzwmsNVAI1qOi4ZOfHuxrzmhOAXS
HBgeRI0MSFyjBSUVSQ8EWwk0NioiVy8O24V3egCbewV8UIiUmixf68Hhm478xhKn
3qqSXfDesZ9LiNdIAl0Sf/IRzqcd3q2fSN1HgdKA9PkbCV+BlUFVppZYvoW1zkKb
+1tHZEV5/VzOmIup6XP9mhCV2JPZLJdjZKYKa4l15T2A3T5zKXfDKY1EMmiCMvwA
VQ0De3EFA9QdSV6/nfBQJB5wPKin2a59YJtVAtkkhgOXaemmFpWsgVCGZEv0JTnj
e9pIMNVF4PwkwumrQdJBYw==
`protect END_PROTECTED
