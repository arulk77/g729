`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bok1EDoIRsFeroqCsP903BOjU4hyaWN8V30Dx4D+mnvGaXHuTzQSeXq+ueLOLdmJ
R3gsuceU2ZMi/wr89UclyVxoEX9leT0Phlfbwr+keKvFA11LZ4RgjaJhtUbXmGxX
qS6tY26wwoceAblxgvIYtB2Zg1uRQnCq8KK8FwNW445LWh2hY2YU5oizHS4nAEEW
`protect END_PROTECTED
