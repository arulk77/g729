`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLeD8VvvHys57sZ3AEHMtm1QfrfNEAuDU61ndmAeGG8o
TtoBSIqhQO2DS8i+Wook9eiXIpYxtn7LtA/T/XpIHbrgO5Mxotv6IekAWjsQdzNN
yTklicQdveGWFVoRwJ8Umukj25WlShSVUfJRRULES7ahQMYJ1pzvt+fDQkh3EzdS
aESRdGixe/FFNdEmCNq0OFSgUmldP/4WC/lHqigMTwxS7V4JNQMiF/JvJtxeAFWQ
kcG381GndFIixlYbqEtGaFL4YZS6CorQHdzlN6MmGnsL2FptkKr01BRt2qgNinaF
iZ+9I5dzKD9pHvChM2PnPw==
`protect END_PROTECTED
