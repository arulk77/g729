`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNYOM1SQezgeCIb+EObLpqWK1MeIfFGCvn1V3zUSHooI
XAZQ1UpUSlF2BvB6c+u4IERhTfEWGLKe2SjihYGtLdHky1DaGKZtZE+WNUd5dE8i
zOLqvNZZmYAEehrQy+AE3O034MN80Aifh0ddC91Izbg1YnNAde6x8Y3ga/wwjlqz
2T0P55MN/eUTVoWtddSH/EYZu6df0HggMOivI6jPIBoOTvZZIUVJO+Vx1rgXsxcz
`protect END_PROTECTED
