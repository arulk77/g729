`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rH8i+zTkJtIuxAQ7L/exbscBczgZ+nAQ/EHvQJaqij1mMwCgnrwU9zNqvYS//uAd
BfpyDuBQNvp5yQZtexLW4+piExElm+1TaKZ4jBeNKQrnzUt26ZkZ3afcZYokXsww
B554JR3D+1ukt96rLamAwGvA8SdEHRefolecl7hQ/wMT4XwLu+ywFsnUAUshkrnf
06JTmBpRWFULs9/930bFGOPYg18jqVBcTxjiUZA73cnkc6PjJleqEsKOr02yOkQf
xZzZBGVkTh4zzcpv164pxjrr/8yDU1HD/L8dXl+qEHWE8b8YFOcTASi50grANYUd
`protect END_PROTECTED
