`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43k7hul63NTlxMh4EiduKvwbpDwWGhzXyLMaVee2ByoT
R9ziWpfrsRQKmaJNDKAOyGA1IZNlLyNUyX+RKmhCqpz5/Nos98vQ8o6tNwGBUiy/
l44nnnx/V4sn1lJWnUNxRYCTljZTWpdD6tU36UIir+OZECcvYd7oTKrHw9s+ZzXI
0ZbNgGRNX5MOziJ+DDNBZXb3+n9DiceLC6njeEsI3CDNljJU0qxGyc3k4KkKWVNr
vaTIz6ulVF/89NInTAo1cnNAvFtugmZX+/WYsl867Ok8e+1XzScxxQDHxICLuUid
6BNKzGrLCUAIu1zhtw4ppwwrSXuGCBgK8OSsQniEIoeNymnMNekKyTbYUN7Xrqr4
RTmHf9ZsB/bHFqyxAfVz6q6h1PG7fQRESMCYzAroEq+J8dmL5G5MRzbY+yNtJXq5
sDbk3h8H/P28tNMwZA9vN4bBezIhdV2YR0qA86BS3mwYCkZwhqGy9qWuyuNWyO1+
UGOMCirBwoyVp0qd8eKqH0MRg3MIr2Y90kRSiR9IS6Y0XnO8+5OSTDMheTNGDT6M
TTYOMl3OdiqOgrM0iionzZhuER62CeUocp+2D2Rq5crQijM1lXM6/tzTD3OZt0Hh
03ouHxTAvU8CBNcLhv6y0xX8KniLTub7oc26DE8tbak37Vzq4AQIVWbcNP5Cl53L
ickKFbcp5z2BYjVvHV6Ov317f55E7sfaattB/pX6njIcqLC2eE3ZUh4aQqbAIlO/
FDyJom8B+OiM7QzGH95OGOKOqZzGBUFdnOXmUsk/DIEOlgqFOxLcKU5EshJbRRmL
IKbmmwwrSueaVCO3/efrDkVXgHJCdZ8QI6r/LPqBfGB5EwyHQBBqXi1OiJbo6z8n
0nAkkj38rTdCpyU/iv83/j4kqp+5UOSI0cNt98CcPa/mIKtWy14esm3Qn6IDcI4Q
0OJ56CpQbsVsFP46ckss6VduGKHd9I0QPRNcc26akv/Dkk6Q3jxX9sDCPoGrsY0G
SZ/Dhm3rPZwKh7F1YOckM9kgTvLgn3vXSKjbcwfnKtdGwJaS++ni/p34KwilPsoP
Ftu4b6pbf0j/ZZXyzGw7+nEL2jJZgutXoZMn3V+hBYwsfSZ3mPZMVQbH4AmYhJpx
nNQUt0rgf2q4dPQqlh0lJ71mOqpHVoRu8xJmwt53s07AKOGClzQRcgXNj2SUMjAj
u2Kesl5UY1fYdUPRI0AY5aCjzrLD4e8sOnTkbeokr9gSIa5j19rPZoUug4OiqA4P
2E9tHrrH1Eu84Km0RXuGgUByTMzMqS2sExg7sRcbdVU+p6/jjIigQ855XPHJAcg+
TJbWFAqskOFEq41Tasx2BJHctQJD33YAnj79029fL0Cs8Pzdd4btTpLfwPJOCFm/
3y4ASYSUww8Wh6ZOw8LU2KinO0Y7U17Gn1MUFw217kfre5rAbIujDrQNyC21vCyQ
FSEpNYwjBfPe6H+Z+vdqrX1VdkKyyxWdWHhvyLAJKOy3NsV8+Gkne40o1lZ9dOiW
4TpF6k8aLKfzqheWrMN6LngrKSIpA6dqmJVZloiX2LLj5KF89OYsRiXxaNIUWXej
ycCHvgmFnfIgd3iIEJV+IMJu3WD0KVV59Af9xLOczgZey1C5gCXdU2IVDnF3kLsK
6/0AZbrUoYu1haavlWUi8kPCUTdQvBBpiAOlLa6xJ9Yf2diPglL5iZJXdVP7NmCm
36E0KyaSPRQAY4RgQL4DMxVO9GiMGRdOeXUjTss1ZEocgYbe0P1rBE5O9LW4MPSm
O9HC7OQrTg6Dkjl3PR84/QGMphMNds+9K/oxb5w/GpKSvzyg9PYFQHwAaMyDYIMY
+aetdVQYiKcA6qmavVpHLYQtj37wEPV6YLyBkSdvoJY/oBZHli/C3aPP1K3QOfHd
0YQguECT3F+8zKIQsKqLCx5reCOQ+Y7SttxCYsU4NM5dAFtaQ2kZ8XwgOIyo3HCc
Q+BFa9LmcysUUd8uaSiwfpcV5CKNLMPqGFDCXTvAYBMzmmn9OnhqJcWS45DJoDP4
d9WGnRV9RR2/M0MSdOpgJi/Uq1ZVEkfk5oW7MC4zWa6tCbFzFO7+jUyUCQBkmCeY
zcW0IR8onep0gsQhINdfkjr8SqEAcxWOuJWpuD3lIScBdY4gPR41qW14eniuvwBk
uqY/w/Wybfaa8tf2AffIbHwNxQ0Co661wKsltCfP+yQBV0uYEFTK/JrPE90T5bGS
Yd+IBO+5f05y5wt0QdOnYQ1RlZvKP/lx4pB0NXmWmHWytOXy+0hfDCznTIqfxRPI
oLmXzegfW5GiziL3BJ13eazBoXysMC8oKxbYvFnqB29XWHuWpoKKQCqu215Gp6TQ
8bWS9tk0ftHCELeTnasBAaQgXWO+/fqSRQvmxqDCmE631/FN1PpQROQ8nL0uaimI
hlEo0kGT22IPjd33octjVxz9cGJx/XPp4Q7neQkj2XeQreMmC7sb+TKgaZnQZcJ0
Cjj/nIAEa2XaOewl7fgnmFP6ykj6uwopP0mRuRsk5vTe+90TKxeMYjXoymCTPu8M
LHpUpOUMafeZK36y3N8hpOdfybwxuzQ1tQV7R1x1ynNP40WBX891OATn6DwWfYxJ
hvp2W2ZeO0gR2H4Bu3aeupgRf3HF1c0tlWWL2BzfWU4p1AJ+cprlUISCeGRHBeON
RbY4kcchxGIOh4J3Fej449vV4cQ/fYlFdFWVZxqMFC+zBfP4A0oiDIoxJzZLQExC
6LF3lXWKKNkDXGINK4TtNG55XvXrYuvG9658FOTxmq9B3e2KHH/WE0BivLSk/JJb
AOgIIzYAyu/yBwaPpXL26051ZTLmVFY0LIEmCacK7llERf1ctCvzCqAj6mUiU61L
Bc0efdAxteWAhG3FtvIIDy/SIEgBvkXDV++x9FKDFvsZi6DMUUhUm8NBvB6xLwKx
d7KM3Bexqxe4jFZFf7fD15X2Jsi+4kpmh0Y/sxMOqxbe5mhb7uOWFAn6ny/ak+YU
nhPlYsTQMvbgliNF+NXko+9xvAjUiM5s9HrczwXTYaujiuW3Kz1u/wz7+i/f41qT
XGrmz+rcu866vNYj4fzApH4TkrrGKF0qx4RBkybPwFP9T1UNN30SSYg0/f86SCPs
1E8EeU9uJxkBBFkwRKxofaN69UnB7PQuD/aEWRppws1TQ6B9V4fmeT8AJSsf3Irg
GHvOADpqFX44U/opXLPH9oLps7LwYOGoCeZTU6hs/xFjURWnKNy4z6u37UxhFmqH
w72xz28Ub4aSEchdI+3auO3/cK5DUA/99xFvd2aWwO+Tj+qhlnEfaOfknPH4qwiC
OQxU5g3iHJxCCTBawyw+EyNoL7ZtbQmgV7vfH8Jx79l0G3SpAPyxNwKQUf0s023G
1RWUoEZNz3Oi/15WpjeHa37kmf2xc+Yk47q/f8MiZG8D2U95BHtD1oLm7x9MpO4Q
L6EPcNi7fZmyq47A3LotTAfG89nzn8WHzDqxn6HeCE8wahgrzsi49YE6o0WKsnRk
rO79AnKYY8VxgPQWI556WTJCuWpLlQhu8OLnfLD+PXIkizMlmktJiAJ8EsektB0y
XbadvlpTJ6tFDcTYgbnXFcy3a12mnX8/y2yt8AG7BiCsWXBOAAstsAVsRfGYpH9X
fPs0ZPa2RgyQhzkFbZhjkIq6DaxaFFkiJ2hc/+Jlnr3uOIN4jP56+SjtjySucTnf
kJ/i5zm/bsTsPoRIKE+amQaUXF75/ZfJfiqW/byF04RxjeOYRzmwVKT3Xr7zFFvI
GorSc1ZMcNCd8rru0kcr0LYbrHvBbCzkJkXpz9mU0VAES3bdRNLNaiwzbJTftMCl
Jt3+cCjABFRBVxQCjth+bECc/68fgUF4g9rki1qNY6VpCkboIWw3pah4VOgJEQuv
y6gbwzOumapeC34R6AkLrD/2UHvtzD3soAcwrLL2WX/eaQTE+4Ycex2OYoE/p9P8
g8bRELbmiDgNlx6GpB+/Of1BlHMjrSiHYgZy7E9sBxqaFdJNejG/Ygg0GR1iie3O
r9TfW8cZAzAB76ov+W7uqRYG43uy2G5tsxkeokhAPTkfUFq3FEFED6ji0H5RDfDu
j2AsW8ux+SbT19XjGF99GjiVxVof9IO71KTd4x4yzUq/5133JcDfTmiyVgO3hLSS
1naZ/osvSqsG1N2ptu6vVB3NNRZcGzoAvDBjPyrsNRXFaWyYYtMZBPyAdFRFVZ5X
WdxM51iavFHPRz1NCEfDXJKTyhRzRuNGJcs008YytauoUhPUmuyXKZX3qrM/qFbI
+0ajF9fOq880ynE31yakynMhJJpv2wliNxyUKD8iJ/ZFuCNK8UnRPjo8TKe9C0RR
9RnZsPDiUjaBpnVDc5SFqTVmVuzofHlqPQ4L/Ia6sk9bBauTG7a+9CVj3QbNh+UP
QlgYoYShiVA7QkShnXrFXWM09YV8qLwGiF7zzICoANDgh8+ycTNfgfgG6D4sZA6Y
qukzGhLXPMP5XUsJC8Ys/4ikexQIavrlPR2PTs7e9KIhdMYvP1uDu5dzbkhnMdAp
qBhT57oUzPu8gS7hdsFj0bjluml1lgL0fP8Nc+bcWFz5ApYy0LNA4ljdwKnupt8F
ZTMWeeGwaU6R6VR0XEbgjaSfdZWEMQRyc+QxkYUeYkjkrBlC8enYBR1YjgxxfFzX
X6q6LppWlzgTtQyY+jl9MFsLydLbHbeozTFA4WppMp80a3PrRXelujoGtFcV/rFs
15JNv/JVyItktMVpR7/8roZ3HrdxSizFiPS4ZBsXXJERVvvUAG+T4QIZoG19yixf
8wm/Ihpcsn2EzcbKeHOmlIRrOB77gVo63y6e1mDHryk8AeCN2kQDeZV7DtPXM0v6
Vv/Jy/3l0ZQ4zQNPs8k4HbofnzY2wNEuWq/mw0JWEhtf/YKkd5T7vhom2/Qxlab/
H1OgYuOKaJeikPzTEdgkSb+EdKUhHic9eW7CngwkHfiXtCJUlnO/SrCNWb/Jnkj8
jz8qfvnY+nR/eqTAxQw8lbwHGI+gf2nhgeO8Aa3H0z+Syfj9pwzcilcofLuemvpq
Lu8RzblAZRcoL+BfXm3tdpA6LeXsnuGItkIrj57Ad1ht6z1XpeWD04SDKJfabuHL
RkuvpcGIji9MZDhHPLbvGjAFrH79xUrwekesrqsFaWN5o4AEuOewn7c5pvHQAjth
K8vecYyOcXcO9V5mMWL6vhWcbvLY1XjLUWnAqGpqz9pB4JeaJnMX/v6RRc+7AlnB
S881GRHFiqtX+v0+mwHtimSxk4ofwu5q3wMAKoguzgF3v0d48uYcM9JT9OFrcwv+
0TG61RkEIM2icR0QATOW7g7fQGtPwxFcnSphMBeFfXo/WiGAfvAYLjCfKmzOF5z5
tBu6rLq53i19Kb6Sph7nmYNVYCx7qhOVGr7rhHbx6Nc5bCzH/GSA5KnlNtRAIR0E
9UlTd6km2zUEpG+DKLB1wWTzwHi8luBLj3loAjgXYy73kle8jxkBEEZzcd3JxrXA
m0odg/COZRiyUH+IUuXaC+F6Ey08O+JkLNOMagrP1Z6W0RrE4G2rBCTrGJNGBHZq
vb4OIZ90t/rU9hZ8SIW10Ki5eE8UAjRHUgEjlddZTp68iYkY9MTFO1TxKpZFq4Jm
FukjkEFNnCq1g/yG5sAE/JN7m5jx/5UWq6YJnGsxqwW8+JkVcqrL7KFvG6hEu6dQ
nmUGaw1iCpFk2epofYw2muq/9Q9DdlUTd4d79/KGdymBxfP5hXrk0jSV+NYuFu07
zlZQVwFAaH/iCy0a/ptxrck0+l4EbL+EWtHmmv4kS5gtw7IVMTqAhJ0VvT6vcHnm
DBdhZ4b+rCT+rOkxBMrwHj+In1zGVYqGslAUSCNPXLQFGKqWerNgd4F4FImbtYgb
I02Oho9Tw38o1GuREYYOgnWyguRXju4SGnElHGm5SrzLoOzDCkDmZAHncW5RK0Rt
H9QvZzB5TMMrNvErCBleBDdnnu52LJPOIVOIESELR2RcnlXxFsylsAiAVGcMb2UE
hP51jSMM49SzpFBgQe0oxJFVOU6QiRbA347f9pKVOwiv/AY+XrxQ1aDHGTXw9rqj
MY6i+aL3WBBol0/Ww0piDPBIwHkIS66GueoGyQCLYRns5kcwRs/FtxFGESjn3Zsy
b3sJ3cgNjsv5/HC0Tyh4A84NeRoWPOl7msuVCz5dIqlEfL8zXbj6B4qJ2u/ftA3x
PheYXnuafrDvK0kMYT+EQuYDeJ72khlWwoqt7oCV0WonO4SFMzs+ERHwhTrfwBWH
lSPmcsruW5kchRSdI3YxqbuPwMKGZWP5Hqyeff2uypP04AGvt+yA7xfaouqWtBDX
pvP01tUDgcy4BbqGSKDhMlz3a4ENUIFQj/RoW97J44aEUqkI8VjoSMQz+U2iACaX
81hG4qwlTLokOLivW7P8rA9MQSwljve5WskCWWkRRtYpWOZP0iQZAzQ+nv7u5H77
ZQ77fSCAgL0WgsfGlxRRHRQjJWfrsO/wSYpk4RcwTGuFvxDfsnqFTS89UZco4xK2
kprruVh5kod4rDOUshvGv3SzrFX1RHz7ZS7ZUa+qKHOXjAPRaSpyI7cGYnKBzOlB
lTyyfkEZyOOnjQaH/SCjD5FAJxR+V3PeVkAHjyS3vNKjDHhIwknrzu6RKHb8bPrJ
eIFcYgov7CZEFrzctG0UqMZQvrUC3XNgzKM8Lu5VqepNuT3hXz7iHHDnDK2moFov
50jgvhUqA6pqPLa5LHMktLnFEPz6/8IJ1przGv1e77lA87CRm3g+Rrv0Q5Hav1Op
ppHuF8dRFj766LVKIJa3oVQB+Y6nZepOF1fujkAzD3bu1HyNM7i+fZ+HH8yQLww0
AZKmjBta/xeE1N+SSRYT/EW8EP4BSMKT3JzuoDiwx2YFtnbUDSXwlHqi96eezqg3
3leS23rV1bJC+awhnRQ371LTOrbqt+HAM+JrYvScm45Zmr18qGh9LMV7j3XYHVJ6
QJiLTYHysgTF0gvc2Au1uvI/PbYA52cxixjSk5TH5m6NYeVdocsqOEucLwth6E3D
YrmVG6fR/DGW55+WqCuQ/mL0/+f/i/dIN2026kUDTBWOgsAxdOfjn26f2KJdAoAo
WhbqnFgeyJc0w7S0UtfSnP6YbaNz74l+OxTmQauiQt0bHdzkhX9yEUMLQjNck+Sl
zhVQieVurmPzWTyshsFDJemO/CI/e57jaT++BkAvIi19qot+cjW09gW6r4KYaC69
`protect END_PROTECTED
