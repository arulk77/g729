`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C4b8ZxgaunENcRne0O7v/UFEdS+zES9UyFMOe7JQI3tn
xsOe+NOD6smTewzsQQjWUnjJNCI6eIx//rCrkkO/TNvz5SR1Qma+fPRRccskcXeb
4lYIsL4vn/be2QsqcmXMgTWOKJlR4OHbSeRSXaomAoEo1s7GKgLF1O7jv55VV8gG
ISX77TFkvJ2ZGX4Z74G00BWSzppGRvFOmNjaecEJ955cJxbcl0QBOOjfFKQgxTEH
lVORiBXvRT2HDGX3sEXi0UKXp0TP2BxpjPLU5gBLTH/Fb69TXkCqgACy44SXIg/y
aRLMgWI0AlQarH7IbpVMaa7qcloYa6msf/Ab3S3raNDf9R3H6iQ5Ep6jyORDFWvY
PzjIn1S+6g+PSxl9y7gwmMBm0b9H5BjdbjwcublFnbsmjOvuMKZfhaVn8nx1a/Of
CVv4KMjTzPv6zZ06YdVp6yVzi7mnIebAk8gHLbCPp2BDEv/32nSPvMMd8PTXzGjK
xsTcEWex6SluzpIybCOQjW3fgqQV+j6jAu7B1YPdIWie2/GsMjgRPlu+CmM0Znmz
L2qi13TGgFr+N3hiIl7sqEYAhgeHTki27fPqFox7F8zgFD/BZ06J6utQ3XkbQojT
qHnHggOOXmIuz8ibM4R1Ls5yNwoE0U8wxbDse62w8zioa50Bl28ltJxsdv8x9VJT
kIQhkoTfqmHqz69AlvVQdedcjb+Gdi363gTiFljrbm4sDtiM5cTxZ783vC5YmpNt
yPvwo42VD/JxQm5VEmfbVmXiQf3KRgfPjITYXMJymKJ2AOY3V5fzHvzRzuVEIw8n
h3k0xyUtvXDcA+I9B2rPxvRIMIEoFg8FstXtMoqzm9kF/rhNKhOG6H+g+lM7bWtZ
H2XU3cdhux7ZhAbaw3b2NaOKgy0S/HkouTIuCJG+8qrtQKyQg1ZKnRW56ncfKfW9
cpeaHynkxWFI87D0mDBRatUijkl17sb2MtC20bhQkrSN3kzWwVHWBz7yEKz1nfoD
ZEUfFfioFJW7uPiaquV4TFmYTFG012P9jrargjOMGLoFgxCYM9bio1Sxspxe1Ead
ov0N7Ii9qaZfKwnLJ7xP88ZL/YZ3OjLgrylpyI7+1u3nmTNmaIv5XbomrlD9cxTL
zCPiIMAaeV88HsQaqbwizY+VdfuQLWt8gJEYLJd2Z36rSjR8zTBycQI6BBfZcUZL
KiXYKd5+1Z76qNEmGOKokH0CSVyq5kV6zR4LI/ANVTjjbr+AU9jWVyZeDAl+suQP
JwmvHgjElqrY5+xehrGwjMMcyoZveIhaXfxcKOPbI7j4wcv+skQMJuE7oMLSIecx
idxA85trYksIoCrR+c5sjZlQh5z1YJ9I+DIcFePY+0uTf64GWL5uupePJgvlKrAR
SUKYqzLk/xie+kWAgIE5Q0nj+Es691bKtIMauY1wQ+OggZu9zGDHvEyBM4tCEISf
BeCrO+awfcvyIjcEPoPNaIPE1E5OgAK6VBY3WKYXHKvLCxUSDssyeLPU7zocBDLN
2FHnyKlPldFYsCUiSq6QxNs/QdKlsyoBjIWJmD/Zs0qpz0taJYz6HOdaxc0VoNvq
vH+AdCrBJRwEfDtEOd6aqTBmXxWO9gp6FZX3q5NoHuk=
`protect END_PROTECTED
