`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJgkoFDsBYWFMRR1QKZhSeJcMXIsGgS2Hid7eO9RsLwv
6+7iVsIu4lc7Q8g/KvO9MIKy/B8AOghKy82PL5/QDvs/Xh/gwg39e38SJgtRlXdW
Ec5ZiofEGcrtlzs+Fsz8yC0Y2iC7MO+Z8johr0Cei1r8fGoYcESpW0KTVsaygcLm
WjpTCQU7BCts52Z+TfxfX8xyN+ugzUonuPHalMq72yDxWKM4Cf1bDzApwo/xZkbY
pQA+S3HCB+fQTYIEv8gUtiaV8dSTD2GIAckOE7hzg/3JSMlU4k7L7FomN/ULfi44
4Mnu3vSIP7G9t45V2F0hfgN9Lz4X2il8hmqy+5yFUCnadC0jntTZqGv9UCLdCx/S
ndERK6iOKR59T4DtSrOVdFlMGj2vlp27s0F3R2shqASlQBorCodwRaA/hJZ8Nu0u
c3z9g7cq8trGvXRvHykDYxgAz+QZXVKycdAKghFC35HQt3SSP3zJKJ9OTgoyg2yy
KlDf9e50NhdLz5/iYX4FDaX72yDE2nk1oBfMf9JbiJDKEVTkR+pjWAjMy4xDeqyZ
h4O98HhBfNU/pNV4p2iQSg==
`protect END_PROTECTED
