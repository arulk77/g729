`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SRiluxZX3iM5qFVgbCTXzagZxol6qOu7I+BECSdT1Aud
C6TU6eEQvN5QA2GYWIG32ixwsUNk+ro6tJTkLSbDJYSWvocbL6vdKZUfCawvfTo1
AN6vJYSwNgAIkzVHaLq5r4+djGt+Xjp0hI6mW8+YFPAt5WCrEoPzpYeeqSJMUA4A
5caa4YWk69H6qgZQ1/HcG0PA5vfu9fSQRyz3NmqaDO+nc6Ul9/ZRLMd3ieIIjNGZ
cvwcWOR6x3SRXsLx/7YBBQxJXfBdGcnhxZZzshAznl3RaoPuZjidFpwU2jtTFtvW
pjwh8zHWV4Cj1lmdZt9nPv4pqLSolcVnEl9VL/AhbVNcgNzkgZ75UZwADXkKyFWj
kY0XKyga766uUsJMJhpGTmohDcjw0Z/AWEGV8nEVgya65PthvW13c1EeR6ICJJs3
apjR2hiWquT5XxQue3pNMGMZSgbZePGYZvnAANGG1SkUCke+sie4Ftc6ZcbBMGqa
kUgnP+LQYpBaTZwy/2r4B6N9z38Clhwd1ARMPwE8ABHUZ/CfdBjxHWNJIBgNE2mR
+vKI1xomBrKGXkju8gpwLr3zJ0kxjHW7skFOmn5SlN2A5EST+BPa5cCdRVpoAnwX
cAWpUL9zcgXF9FZ2zBMFR1/+SdeTp+f6E4i5B5nzSwO5TKkD/yrDKEoGRV6BZxpn
MTPokZ7eBYm1D2tiHO/SJfnvKi3UjEhdvGRsgVUKPf+rgKI8JhgzJpc8jd+Q6j9b
nhx0+iEM/rxUdGVYPu2nKjB6QB83kkJCsZY6wEUXILLEXofDv58bIh6Vc5PQfrM3
bWVG5e3qSsImu3OEF5Z05iSx/AwfU7ZwSGdBZ1CE1b7hUQrNscFocKVs52iP7iPS
Fg7fxzeQeUrAeJNDqCKQTbru3zF/tutqm/RTdX+tRZMsJovLmSu8I+jGrR4u2Wuc
DZczZSWrtcet0nRblYKaFxeKBb8wLRo+Z62a9HN+ZxWRrKRyGCDR+IfVuhZXqrN7
7TMzanWhKZi8IQcB72tl7A5YXMPu/SYU40hBvKcRQZ5cyOQbZZYezLtpvLqzqLq6
UTBTmI2xZREhhXKI4UHXzOLlzVlV5ZQKFtBrF7YNqwLAodjbPM7qNTvdunKlIQeC
Rq+fg7PQtU6QPCZ0nt7oLDzIQ8EBtyVPlJZqzSD6z6swf4ajMBttKGNoiDnm4lS+
CF7WVcY6LpMc/1afGYG04VQk0o4KMadRKrDglb7djOJhnsvvk65HjYAtRWomuiWF
BuBqjkQtZkfUuP29ZYsjqd/V+Lkm5ubcSxvL/+DHeEamwI3RBiNNLwItZOx5l5oU
4I0YXGdblzb21Tadz6cZ3RcSuJ8lYs4tUUNuIkUttD/p0PiSCfdpeY4doeCCMk5w
V2y5Y4T1TTVC4icXN+lAFDA6klqjs8sGJomqZjrhvQfcXxjqstmJtQICp+F4udfP
lI5/oApB5WB5VHAD8d45KBaQ0sGCH8eee49G4rsEMPoGR8plmsgQHJzgpMUMkt3n
w7NVbzs/od7wQG5oI/3B3bLuZH/4egtQoIoFPxsFtyjg8eqrC771oyt/LAWKOme9
C/WtT+FoN70K4dtQVfp3C00ClGW97TvgHRxyDb6wFhPid4ewZeSmd8mjCMtBbhkD
K5LH1jEH7/Sao5Fvr6zNvgnmCVbgcv+aVB7yv3HFzcYbsqEYY+FEUIb3+K1IO3tE
6GGl+FcM/1vEXGUWJpD52cYERuwJgWIPAEwZzraUP78nlDSCURmCt1mTdXS/FkVB
IzQs+OU6w2TpV9WaCeJvNA0kcGzlAKnEDPKgeG+QYEQ6dJGyQlR8OCwwoxRHPDy6
SB52dvmDZeMdf9f3BW8LgrM9dNXJlqeRyczHahiQB+E9o34q3g9+Owvta1QVXA+2
m7Z5ROi8s7AJ1QCYjQCnmV9+2ei4jHHcHdrJOgNS+b3fsVXeMw4W3JpP9XXwboKX
r6sfV0rWm5SZPuzC3mm7/BjuY27hJ7jXFlLNjwbtu6aWg+FrlWnuiEdBE547jvB4
Z4W19LUbCNQwJy3NftOftpMhWfw7Aybx//o9q4To8Asdmt1b4bcaalupKsUC9Nup
I2qXdL1Q5rJggZHFKOB5mhI/76UZIH9rz9FaQoABbo1tn/ybz1fYSyUuJevpOUlc
vd/0wqM5TV7+wI/eqKV73s5uaPGIZ+d4hvHU7298knU4QcgmbA4smUtme8pxM3eS
WkTmCl3IwcrPdlGgobhlkO+97zJ9qkaVSPkt2vuU0Wt64ldqLwEjvRdAI6Lo4L2S
Apbh7nM11Nfxcr7lZc9AkS/2nm93ib3XeqqtDX/+jpPTISXVdVWioL/kp7BEe+DS
wV+e0wUywqBjUib4bgVXKfcxnOEQvmAvTkBr4Oqh4iKNXSOfgnWXN8M0MFn2E1B/
IHmR28Ax/L7CsJ1fQuI1LU96B9zQ1D42ezeStLRMAfs9uAdqCBqjbwH+iJzuMXQt
RDi+OVWwFMYy8diW06StWB1bOpaQRf5bTiLwq1wj8H56MKuujN1zOKnKPPP13/Do
w+BsXjl9FZYRCR9epLZA4pC749Gh8gfmaE+XvVyaMKkLW2fVFqtdK7K/r4/GkhrZ
1tCZ0ZvlsxW27mf/FLQbicq1odFk+Nf2pLG8drinJyJylwgWmbDmakD8IbwvGaF1
emXVEtU5yRv47RDMrc8ctwd9cWaSSxGyzBGDcNC0xoOWsqNYBD4VevYgFPsnAsAi
HHdw3iiJfwcCJjdD8MqaCR144YlxOF1KRdKAGcHeBxKoRSIGpsYQeDhjO2zjKj6a
aVencOcSha1Eln8+bCtA3en692Lo2CBm+2KpQPu5GJKLniT8XgS/z9D8RY/T0naI
eEsDDt8bV+poOjjkTgjdGXxhI4JdKw4Iu3tKfskrb1r/BSlydDASapRoBKqFfBEU
t4L0bPgTyZ5DDnkiY2OIzwR+5l1Wm845CCjGoKOxBX8ok6LA1l1qeOZ6kTZd/QHy
xPVDKxUHG4fArDkOdljr70HswuufzGrOnyk0TqVIkN5dilRDUz2hP09gp8ZH8qbJ
qOPDQk6VDzNtT1rCpPgeUmLCCJr/qmosp1MVs3YUpFts0lRYzUu9ys3kN8sxZy/+
HQf9l9fzPJcGBuUucnzToXiB3V7Q5HRAjl3h+tIhHO5Zv0JqA38bqoKZc2VStKhQ
PE/QRDqaHqz64BD/szCy2/FwlLYzdgrVblzTkJpaZwstHmTQqpL8M6epw0TD1NVD
t4C44YN05vHPU9Wlk88Vmya2ismGZIEqpIROeC21qCyPkNHMad2/ThjT7DqB2rFB
NndbGs97k/+yxFAGb7phsDTeF8KSku69ThCr81WobX/trFVAtsjrGIGIMIqlBnPz
1uK2rfBa5D7z1KV96nEAhxzd1fJikelCwjwgrZVohS1I56e5GggFhDmofRXfWaRe
eCovq+uJKvwdBVrsUKTqEeET3EQD4ocO8k79OccQlqQXHE8QbDIm/PmSM9ri2/nk
M+Iu4Xpdw6kl7kVrxvDwBaYc0GJlhKR8J2kbtluXi2h00Fmc2CotdOeUL6Z0E4El
EDYfHjc2A2l+HfFPGduiH4Lu6LNQT+yv3AsthfpKQTzIyqSQH5eIwcqlO27VcYBV
WNCFLQEf5ZC1tezQu3MuEAFlWuD751rGpFegE2wpGdCRkbrmenoCl7C8Jn4855cf
+2MbbZE91/Ylqcq8De5cPxuP+wOb8E5a+d0lvDFzFHw1uZ6kSmwaKyxqZT19mFLO
zOtGKZX2rXEbacHdiwMyLK97ol//kT9V3g3MZZiM2S10FNQEyuQW5kEbrAfGOUE6
Po0rY/jCL1aScLXEp5NWMqkDKkJaZbzpg4IWH36mGnAA4x0ur9z6uG76VXdrjels
O9KW/0JwnO6As5YvTXmEwGsZpiLTRM04yZXKDnAlM3r6RF8HykDkYtUoYGqNfyjw
hwVzO0wc9OSgJja1iugfIjDDQDoiKgbAcNfn7ljf8XAsZBuH86A8y7Sq0QIEFH+w
O5w2BbG9GFzKkUWSXPeuCUwYAmo5WLsKtjmMZ9WeYHdqmje8UmKhG0geJDUTAfzy
mirkQncbKBIIrrAzHTXqC/dlCOytA9BlJNuFaNDKBirPLJD6XHBDx+HfyS/WtEmT
lTDiLDhB0gFGrYbXn0Q8D5DeHU2ViysoJ8Y3Emm9y+afIrOOUeTGAGpsqjRNoTue
SB4Tto9i1bj90wl3iTh8ZZACCST0UL2D3iTMYeHoGTPM7tm0IrCN5lTs9O5IU0kJ
QCqOz5ubhp6USHDzntkgkxEogpvd9GAObTEAlJyzbsb6oQ6TVpjp5Lmp9Qed6Qru
cd3WJoKEWL22l2tq6Y4l90qnLTRySe16ULopfn//U51b3FKtvDllXf8vuqWPyThE
ieDMPpTwHQKYI7Uqz64+WfIhdpKMCmiKRiybAqFLqYoEFX7U25Yfkd7WcZybV890
pJEPFE2zrQAYW2p0Nkggkq1MgvfK+ug10068aBylXEXv/LiqEd2O7vsAJkPI/lkk
fBrXM5AWAX50V7GgRWc/vTld56mq6vN38H9OzrgUZl+kbN2rDeg0pzdRj05ZtLN8
y9L1pF2p/RiIvcg6whB4lBTAiOUtPitJmwSNHhiLWGyL2kiftEEqNo46tNh/Nt87
GogfSJo6Cx8RHJNmzYNDyhaGrEYyUTM82sTlthXydJdlIx8jpRfbztRlZjYuRynJ
PNu71B38L8rDCjqKGg4FsBXAtgExvrKRYOR9BkUr+GNJSCyNdkmHMfc4B8hVyD+9
IHdZ9ShyBE68PDTuffLTyIr4jHBiMyCgz1h6Tu3w3FnbK4QVZlNslttl/40CnyKk
jsGmhtltZwxlMENApi+4lVHqkFI16YJVD0EHFf9HVTVNiKtK+xPsqvr8caiGxWDx
tSQovEJ0E5Xq8XJDVfxHbO1tL0qXkKkhcflV81PCZ54SfDlGiQCuEs4lB6aNzmWH
1exdweBlG2rRc+apY8B/2o2JwB0xZsjkVwE+aN23/e5IqJXojgcKqZXFORQMZzvf
AUc94aa/E9AloJhGCgZ3OasK7pxOXku/ZZ2BK8w5HaFAyHM5Mu//TMysoaQHiHtt
uY51gP0sCRNA/lcVZ6Er3pU7obv4GB13V6sDLIMnNwH1/5sfAMT3piDQ8EVtcGwT
4LneNRzvNYHsEq2Kt7qGrwiHm5RvGxpoXhffwXZ0uLiaLWsADw13Zn563j9BRVL0
xo6F3QTpJ7pWovhLm7il3FFj58lR3gWt+qD6LlTWYehmc/l/bNURLQFvtg+Xt0rh
8VMsvnyxZ7kYpiSMsZ2dw4BN5OCloSMs5jaX0pE9q71mOG/xb854klVSIi96H0kO
+XOWDlX0gP7CnHbRrRRmyL41wXPgToZQ0x1GYNBRIyM1uuTGk5a6zJHpLX+KKDdh
9m0Q/azyvIp4LZ1rTs2mVDmcpTwDtYwBobQK4oQcaUHxBpwrPtZWpckaLQ9kZR1E
eV0Gkn98PJwePp2jok0I7RINaZowo8l+jz2rE2Q5D2eaWi7f5aNKa4gTIqVajhi3
J8Crflwmpo7vjrCvh420HoXI81pjjtKN0bxa8/gprGMyAiaHSBSOFbPnIcyyd/Ut
hNEZ22VGZWshhOt00UK64+LqxRz4ixhhUVj1p53jK5OcpXZGvz7zKTYAu16AeBLc
QEkPqtSbrjyWEAHnf/gnYMHSSlBnjSkTkWsjn3tmjdWawjMybv5mXFoFq7uYLL/T
jyQ9HMR0JUYqe3tYgUL3hSAHb4SBetw9RzJNXn5QCYTodGNk76PMye/vMGKdCnlv
fzne49DMb5pqrosPZ/XjAROITliUfkQuncu6IkkjCGnD1Vk4ORlyN8/oqGKNbd8a
N1OkWmGQ+hCdzoh+A8wKheJp9BztPIfZiyIiTYs1FHKDL7DO+V0vnXE79SzKAFpl
gIL1KnOef09vqMECmUUZ5d6lDtrZaXQ2L4P0aRqMBj+Ze9w9z1kJe57YpJEDDMUa
2eM1tUyKgv+egt1F5NLbTlwlzDb8s+FvbiuTvic9AbFyteg/QHm2+z8wOPm5mzCo
Akw26g2FL7ykjQb9uOSDJW5Q8/Y1HZr/x8pngIh712XXvtW+tjS2xAoxfXB2dARl
MQD66UgX/OJtsmodSlWydk87QwKJ3GauTIiyahE7AHYvmI994yn66wfEI4UinLlF
rp1PDR1ri3glUmiaO3tP+sUpJ/rCQm/TKWd/akWZJcBPoqX7OOwf2J3VxenrNnvC
+0NwSUW7ROpaIHEkBaXw+u4CAJvAydIv/VMPinzp1TwtM1Dzk1EIY3wAkGqVb1ii
/QcfKo6HjP/CVLUfHjZXibZTs4BQScaI2Fyf0ZVjTaZw7CeaJu1Osq8f5n5jvNuN
WeaBzHfVkCd4QaF9uEyLes5EnCRbrUo3loGDRokSirTkf+HhaXABpuH83zPJYw06
jaC1GdnYRki1thrj+phKQxErFcWcyVt03LJVsdeIQIng7ngRyTXMlqOulMN69m9d
eSpmFlbxFUbceTKDEMQNN6pUzEpwT2JQPlQFyVoqZt7oAIoVo/DcrejImXOAVip8
bqpMaGSO4yuYPbRO6uLhZHbv2ACqaRLDyAj+zqLp7UzV/u4WYD3OZ0gLZg5VMaZg
L4WypHCtvWE0yOiAIEC61HDimndzRDIshC+ge1FohaAfEwobt3gc0EfjMCOUOOKG
Fc5GCFvcTOm1buH1MWOS14ZXlSe9xxK883VhdDK1fifMs+4ikC5GW23ncWD1A+ek
EzMhB8zaicgPwJ8kjUakuiYp0+IJ1CflGEk/XSvpfVbM16nTkMo2ysi9lFDCPMvu
vB8tXa1SXA7QnD1KByjjecdp2WexzFHy0xIq9mwSmpHSVzwcp5bF4U4pP0fpkhJN
r0mLdzedewbSRISmukz+6ky9v+YsudkRu45yQKpJfrRHV545KoAlo9IF7iOZ3Uex
VpNsCHPok30YK0/Ut20Gh6vlJmAdByYzMpCWaog/FEE9a+T+jwfGwuX8jt3hX8tr
JbzlI1VZksViY5yAwtNjgKf4CAyzNachFnsjnn1/LqVqnfXKE+PzWmUIHnmX5ta1
oESybk4G1VmvUcsd86cjIwR63maM4xmcmB6WO9GptLCXRqItwMpBG2TJ7+Q8s+Xf
P0cnAc046XM0JgF04G/Zy+ILXBJlIyLN0Qxmx4tTHsZvnHLpHXJ3z1OFZe3d07/O
K+P1McRHGpauM4qt56Bz/fsySIvHoFmJL3i3J2n3WP/ZrTMrMt/cWo0i69/CEOTw
KWec5vpw72AgIY93urC+xwzHxkWhfXA3ifXkldDjAUuBIiKI+jgqslC/sOFqBiit
vnCQH8bQeEs6c9xaV8meYaKUV5ig4mTynSGw45tHFPWtm9UYELjrMrGM1nJzaxKv
fM82a1qPWUOtu4hVnJjdoRosmjWLxu2pAY7Ombmqp6ijTCVB3IXd+Tk+6fursJKD
SsQe0BmRCRlFL49oI7eaUPCr1i3c2aONHbnneQ6t7KYv/39nw8MCo3JOgJkw/koB
zFOgZTEKp0oXIDdtynyq+fnwH1cwWxmenEcPziLPFb+fLhMyiCf3CCLw9h55suBA
k29I6JIEVh/roLRJTggrQ4b/6XSED3+fyJ6hrdA9QPTa47dWT8vnR5bOoi+r3DAQ
k20TSohxogxK3oIwUm9QRGUqGo6KQX/+j0TLiciwQLd5rQOcnR6f3aL9+O4UGVFB
qJTKf0HGKKBMn3rlOM0iJ4QTAb3rkOFbwnMBsbbq3gHksB17E6J9sJcNveFVITZK
U8mR5rqqx1gpik0epQE2dRZyHWlrNvC4e7fVEBjG9LjKJNxU1bgJ5vRCmrn8bdQa
aNrc875NbI1ZIu1ukPqeIvS8XkUGFuKqB0xkflLfIB/E4cyr5jrsB0wGnaDyG0Yu
vXgZAXd8gGKUoJYMCsevuFF55O22mBW5mxSqWKMDQNMDSJZozcOAzKqQqMicFh3f
+9WOzc4CzxgDyTUyf89Xk5T5L2ZU5rk+OzlxyxC6TgDq3A4gAYL8PJNS9droIeH4
ImlMUKkJgHdRd0UFpQ/l22GpHtcGGqyGv6t8gD+s1lNMO5rsrv6YL+ske8u/sCwa
hXab1WWs0pSW2sSyyTuGFaLI6ys+xQdmXia7y3VX1mA8OHMBNB4Q7w9fSTHE41Ia
+frwViiYf1WC2Ye2lSS6QhkQWT3RkDncPa11wKI+T6znrNaSi6KDsVqy9VOhPsP1
ueNQBGZj7JN61SKl9OsO4SlCTttsuSEQIh9TOArBhpo2DtJnprMZ+79AWx4fUg34
oI5pKPsK/HhT6oLtdx0AJdaVPqwv7+UT2BluLkr9Pdnpeu+C6cWTvpWEZa0FK7zx
8h60/7skEsjRKmVUNazSn/CnFvpR7ruFtpnSIGBmYQcfOMvHkBss+vQYMidJwN4Z
lwBjY6MC/84WmYTaLvgWx2X1OY1TcaVKZ/vK/MpOu5fFDew2N9nbMv+hV3UoBLSM
vAGlXKM4drsNGXg8qvL7c48WYARAuVc6b88/Xoa7emhW4pSh5RFQ6sBDIuRWU0dB
nWJaEcYAlrjDhGhzCu6jW77r5uo1F7BdyinYVrKgi97IFXqQsGIz3/yCMSookUaU
9tw54po9csgB6tl/3IdNUNQtMv0jRpY/HU98NJl6mES22V80jQqGXp2reqrIJnwz
OW0H+aGkvKZHTrnOKFGiUqX5CoiVfpjr7FuaqMBq8qSVkjzGoOwgouCsQQRMjig6
G/rvY6CfoDrMVkdEYo3rpJHdrXq3tcE9RyN5z5QWctFP9pBVDyhWvBjQL+cbbCWK
mbK1lSjjnwqaD1DyGZr5T77Rl/gX8iVw2dZSrirb3uKA0oa37umR9v5iXRFm4OkT
3UG8sCQtQIk+HmmlLjMWtD3rW8PjJW2kwgDbbsxkvT5wQDVVxra6EjFTGQHg+CmS
sjLbMsgjX9FGO3OkojcpP8RRar6xEsnNOh49NQb7vWR2oVKBsixalOZGfmsOXPfL
XkrAc4sdH59ykI4++H2A7cOnUuogcvwI6Z3rYuZzuq21AC8oblsL7o18jSHJlQ1s
5qRFtj/TXuPwwO9AqlCycbbkdkKeUZ1EBxAHafZtTaGKx/7mCFkOOCBoPENRtF/H
AJ5jar5+AcnxaWb9GgMqd/7x9Cx71xcbtMD+epolMNkHn9M1zOMyf0hZFPeFWYfj
q0OLqD1lVXoK3g9V3qjN5324doTF0LZ6ZLhUGEEDgdMwdQPdaSLyXtjvxSxYfmOS
cdsHzWTD0oKQ7rDNgLwYPTIUKuHY/BK4BwmsmYSu3jCREKDLoDYhpTGi9ePDk6oS
7ABa0TZp1YUfBduCV+2LaUBlpDWjDACBvvCwXL2f7KNy6W19PdIsz0+KCqEicrwP
/F1XQ+wUCz/kLj2Hs1X+cgrq4I6iQ5JYhJS4UQINB5j3kJfESyjcu1VblRD4B+0J
tBGzOel8okf4x+hdmFvsoPfgW+PSrloE+N0i3CGeSfp6xb32k+PdJ42SbABZO6G0
HsLG5w9ZCiye9XI6ZPsGU5MlCZnBlFZOQ0U8ACxb9ODOcZSlSnBXP7cPyK6ptoSk
uwCDKOQYUG29Ad2u4w2tIw2aUqxxtaOjbJ1srq2+msbpIk4cl1yATLiTI53baA5x
ak/DkgXIpuZTulyKi5ePGXEW+bAIiakyoMtDSv0eZO8Q6KmxTSfsjQtagphYIt+3
0A8l0HfoWt4KCqIRZ4Z9VuhEfqfjj+qaLOGayQMPf0nYxOuIcBPisMOgJhdDXS1I
UNf08bZi5taX57phQa7ppAE+XTfhbIzz+3c6ziOJGIifoZ3WwY1mHRqzou4OELZ6
VFV0n4I72QtBu2YdGW0kCv85MjR/Wb23QDbJt0eX9AlpvsnDe3TDU2xklZDf/hxc
m+ND5uaQNUnl2BYZLAWHBWrezxFLjOedVRZoAC58HLeN3g9aZkAIukyWA/DEqk9V
ugdmIVr5srK9qB4ehQl4rK0723misH0aYfjA4Hzxm48OUkoojL83xdC5YN1lrS9r
DX2FKrYURAALFv8PcWSzmv4w1vNaX0YtDm+C889qersxlnA0NkkS+42trcSC7dQ0
uDFJ7omqAvdJQxNa/G4O4k8erDpAwxUwZJPgE8mFpYc3FI5a5YTsbixj/hGONeU9
gl7jNW6kWVfOFgxIpbdbUOVHw+5VKAksjqXI9LJ+Ttj4XKM3CH1eb2WjJSjcR883
0P023H8UdeIJc2MY8ykG/CGb98UPfK5z7VoPOPQytzjYL7DqlwIBYXru+flMRmNb
qLLTvxS+uTcfNYFdFvANUBB30V3wUPu+keCxRfXbAWgGslZeXinpnD0oDo0G4+Nw
eiLKNc6qKGol20md55YmN4WJs0WHTBh8Vxml3s2XYcBfuRJSDgjS03kSHSQpxGiU
uJVE83HuKSb8N/hjvAJVtlJtVnjEa0kjT1g2+Kdsgt3KDYK8+FevhJI1IYcZVgl7
uL78nsuBxiJZQozhCWFOuBa7omyDOwF48Lg4LY7MevWyC2+cNeJ+jYiRZg4nuHhi
+nHtSbyVK1AmCCprTlEwXwWtTD63H8tmNWOr0l5xJVwF0xsS75+qlKN59E8gAyEB
ID8b/eNGI84Bx4GokJhhqXuLMBIdxsNYQPnyAxJbFPJ27Shkzqegw37geQQBOw6J
wVxfTAkHpLW59sRdSzTWZcITSSOi0kemKuj28rTucW9XDhLASvtDseVVgAa9z6LY
Q2o+SKm//xVesLyYEdiDfCgBfYeirxdRc0Cg14pT3/mNqWHH46/uSE2Tel5M21gi
Xj0UvH9leiacvK6VusU79vEOcRVInq1M6QdltOMul/rEC/12JMwPjDwpXoFR9PNO
ypgLhAwok7z73IYgi+O0nweK/Ue7TGSgcS8DDqrEBFVVKjGQpoTwYmFqQSlG16jM
WEoEawYR8bhxiAkCjr4Q0Gn6KdVujmyM31Z6QK/eJGdXAit2AKQbK5lXEwb4PzbE
zzCUT0pT+6ynlFdHg8bI0FLgEb3Sa+ZGLWHJMmUbjsiqpUmbS3geLk6m6HqxlKdk
ozJPf/q3DTzg+XvCGjQcsBhTxQE/XFTOXfQyEs48U46I2YHVqFCLWblkaLoT+lF8
YA3vBs5o6ZHy5OV8yskn0e5hIrr9IEI/0RQOp/UIKW+U6RAHDydrd3QQz9FshvZz
eEALrAWBNzCx5jp36SDBF5D0mC0oIEGD30ewRzv5yiqouRUdTsIa56qczC31ZtrI
qW2AkewQ0h18qoEqsk5mlyDpCNfEBOrTd5J8FxHyM+GTEdoS2CnKA3iM+CvIHSNk
pOLmE+QxbjKj3S47JxH4/ht5b2O942R1xpJ76KCH4HbG9S5gkTbrC479u1JqRtvW
vFwHGiQzo+0jne6i/XZb82UpW5FW/kowEWXRaamu40PeTqO9gCumR7lLB/TOEi6j
UQqjA7AzXmH3tWRZ8ARhYNiDiofYFlvM6fST0+OUbeeP90wzO6rZFcUdSBAFnwLR
JtqcV7OTtK0GeEh4EXcuE3NtNGZCxAoIePinuWDZzEP2uiaa5/6Lzi7co/bJk55J
9B9sqdYYpW827IQaj7f+NWFrCTkaC60c3Y7YLK1MZTYqhj6vS+1sLfxjbMSOGj+I
DfAZfHnsiF7ku3amVWRWnxtzCF2T7LxJ8WDnZklUH/ACUrMJsBANIu0ALvloPC2A
7bpuBssIQnUWJiARkdxkxoLFm5uzCvxuKCnnzxNBrZbkPCYmDMjPKmLWQa9Jp+13
vOR5tJNMzojdPGytvOzaNM96lkamn6IdyokowKz60JFczaIthb0PJAOxFh9mcuYQ
pHzNYkyfPGyTc+FAOtcSfB2D1VPExkYuHIJAmBBkkA8DVoJxt5mp+rD+AP66q4+d
h3DFjrW1mRqbOrTW8ewXYcG4fAcOwASCDr73g4aBSgb9FfhbmIxUWH/H8o/vfPv0
F/CNgf8nelHTuNqdDGQnZb6UZFWV0h43jsGdImSo3YndkHc1CuuLssXU5Rp3iEgL
TtKKie12pyylnCZU4UCcDd/Q51UonDqVhcRc5yqlm2loVCqgCYtoZlnyttR2rrMk
16e29BYRUm/Sc9o0hZ4HAzdFXf3kPiQ/Q78KhU7nJlRje9Gy87Gm1cWk/Rs8dQZ6
4AmM56kAe1osldrJCP4ru6uvhnqY9iBEdwGpJNeUIcymnx3UMyhPGVjd3LDLpwkz
nE24ss5cetIZIw3vZWssW5tass2AmnEsprtRCVOuwJsHmRS7ZYq74FbX/VPgvPhR
bZLfTfmKBDZ1CKap2u9KyjDVJR85IZP5VJvFUMVEWq/J+hn5PmnqpmZF4pjDNPrp
2l9iODLx71YD/iju8qSZ98CPNffzIAGcHpaR9R9hZcdECp3HvwF8FP4MD4IvGZdb
S68syrxJ0TnlRDZLA6H5ENFB00K094w39PTaEC/yElsgMhDRcjHNUQi9H6RMTBBc
dJfN5vm/GBvQz8lBIH105Q==
`protect END_PROTECTED
