`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJie+aVhBUd6+raUsPHsv8uUVwN/360Lnfoddse7j2KA
CQX0IGauDPRGXrEFgbxEe7hDhn90QZoAOmU+sVD0iN5Ruy+j1pwcgzeE63Z1tAxH
vvgFZ0rFDT7ubq4Mu4Rq90mc8dcCLGfmtFJiFNNEV7YzNj6t7RwNAfwqpnpWMl2f
fu5aGvbkgiMCwX0v3HJLf/AtkC3rksdgmdgXS6QP4WZDezBkHj6OquP/VqWe5oWu
UmCTKUbKioGR8M1eB15R7bFa9+2skwznEr2gtoZtwB+5SLh8RiwX3EkSTaY7CeG+
n4nSEhlxHxbiYUSY5HWVgUmEc+LqIr5W8Lsv81uzdNattD9vt1O1UdJOdnfeWTQn
zvCG46OnyAFjMAjANJ2q2mRKWW72QC2AJTgjoRpY8+87oxZqGIuT4psR+q1d2GIu
BRk5MvW6HByW55GrbstqB7lQIbUYW13RNFsPxD5SDLJ6DghcLjWuaKU/1mMJUgiQ
xVWsApz6QqGW6THv9JR4DOvSMigncLr53j+ZuhMzqFpuoM3DyEeCdZu0/LHWG0Lz
pZoYJeU9zoCVPudrmIsp3Mmcw1mVbJemCrO7NU69JcsNnJBvEW428IKzUnhIOzkr
`protect END_PROTECTED
