`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME91DPF7Zj5NFgMNBDZx0r7ZRmxa/5YkK5AhJBXwo2Tn5B
amvXByU0Kh85qiw1rrTOSfZTLp0qjfQ7SMKCffoeGS0K2EuRt8goAIm+bIW7z9+E
NyoPwdyPc0DIZosSxnMI2gP380aJk8BUEW3zXRYQYd0u/OSwCPz7oPqZReO1+ZJv
EiknoL/73bWZhPdaKLN3i58/f4egxKUagW++GZy4/4HjH6sgYmbkI2ik0gYFHt+/
UfOneWKs/jwhzdqCzPRWuaxaN5QL9o+IZitBUKcsb6bYwJxljakrgLH2Hm8zf0f+
`protect END_PROTECTED
