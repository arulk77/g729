`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMIWUBr/HnTzoKeC0MkRrrdQsDVzHzY/BrTevl5yZ568
ON+KGtcAvGzTAE3qBm3ps9vNahGDeNR02K6CGGfbcJg443k9b9HF9SA7mWnalo2q
x1oGYGwNnrkxZde/uUd2aYrY6uHYuG0uMJJEO+4Q2mMsSAA/MWkaw17hqXCDUUyn
mykcrW09aTUCpPyplkuukf45p9aW4oCVNEAK3oGXMUL1z5g08gJXWNUSrsz/0589
ezqqmildCqluVLHhZO0NO4+Scn49OTsZyomptnQ8+/d4agGP+aUCUxBRHL1+oDBX
Fo4EPP+KNga84fPub/G8DirHzLRYSCb0J0uo1SdkEZZkDeGuXoe5oGwlESjlnjQv
nGzs4fPmhlSPfmYbVpYzPxDMZ8yxtoxrzZB8m1OjoHQQ5h+QInzWphAoLZLsANds
HdCUcY8EKP8H1P/4BbLToaoqybuOlag/zCaztA/15/rm5eoNONqgwiCZlyf3mgYC
IkVWMXd3gwWJWKamx2529/wg2YbymkekWoDp3NNKheIaPVPcDUXBnFU0i9tRAq11
BG5tGI5yEo9tasKrtgJONMqeAjvo/++qLe9LBFnwvb3fwTN16NVfDKp4xsIJe+2C
yIggwqpoaHH7PCawvqRPtQcNVPEk18hDNaPlBYBsnnmGVORO5yHFgoTL8pTTY1RI
3uZv/i0ZaS44BOc0J3vRRZyGYkgzd32s6UjK55LekMGc+3kT1HE8SR5DY5vM8zoN
Z9Fac93WK/tsSIv9s80qr3Tq830EP9/cFNXeZZBWfSzS7MhnyrpbLzUG0yccQWIv
jJxtl7qQfYB/DSY/XO7tldoTFStFoc69Cpa7cFlpPZuvo9FfyuKbr41+wyy7kB//
TyNcbWnx6bgnpnjaTo0Y6kIsidBtZUmh67XhHUgvIbV5Vq8Uyigp/SFUs3tJ+gj6
`protect END_PROTECTED
