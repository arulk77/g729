`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNDC4r44i+57GVTqkFwNukhYpg0jCCh6BfTn6NOeRx9p
HZntMmsR/6C1D+knnmn885yEqT8421EpHfwIXnr4xwm2dgz3Xb/FUWDsYjTVg9oW
RcE6NQpWKvd5znTLx1W6dwELJm8gAPHPIfCK1s7l+3HDYyb/Or4LCpcA3udc7Zif
IkIST9LIftZe0h2cG1ULtYyghdDDQfjUmVPccM0KOULnxec1eX5/pbCm7PX6eZwG
S3lKCCv+hamMHvM87XKhaX0ImkkgW6tuYdew0GoFb8TcMMevKoa0rioEPhWKDYfo
p36K2ckLF0fs2KrmfyeccBFGf6cFAohrTjc76J6xsFdENZ/PoUufHF14CCpZq99T
XzM4CX24yUsyNHOHYCxXm08zrus8W1V6o4eZ9DmZPNXqJvWqyxrx2Fy9YlMb4Z2h
nICfyvLm/ykEfMJvZYhVAWUsK5guTSHQBjIRf1VoqpTG6Ccz+VPQ24f0OmKIJ5kc
hWzoxMApONCIgvcMhvJURV01mxOw2M09jjrnQXP+JGCq9i9Q1rqGLM7BKi70rEDX
yj0bvjl0S/1+RxftlyfNCg==
`protect END_PROTECTED
