`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wJzsokOQhWbfTsAQbDjgC9PoIEZiTjyOr/AythyZFWj
91aCfsvFbpYVQLUS7zQW0j3JOZU+mtMH/MVH8OMJaBbTs2YpufvDB/uuFf0AaBbN
KFm4dD32kW8gXnSzMoqLiuR3S6zPGe9TT4/zVDo0ulYxmeS5KfU40JzQsFrxIVNe
d0Z4GH4x4+aaoiSZRmFgeaPmjFObw4Heie4iLt1auldYsebucDCLxbDeKpui7MhB
9VCLdLouXJ2l3w9vcMMnq+ACj9WFh9l5CDRKVwC7nRucwhFhg+Ouo1YYkeNb0OCo
0ujp6gVDudM/gNyWHZu5zQr8I/jOF38QH38j6nf6s6LU6ZAeXLuWx68brygeB5zx
o3hDEAe5bp4J1D3OCBUXPw==
`protect END_PROTECTED
