`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFmTNZPM0+qoVa4U2my6eYlXpT0+zBojcdpt9biZ2oaY
opEltR0oht6A7O2ISDxFzWwQxFdJxVMufUu0zz+68QvpPzY3HTpuRKS3MumhBfT7
ANkXlN38UE+e3uUl3lrvCzLmvXBlKp1NvkvHGY2YniRYg6NwmuvViT+vtCX6pgdc
VnIQ0o4lxp14gOzjtyyniwYmjm0/UiQCWniMDwD261EeOgsvZGRQNW5oYgXOqRWG
FsMrAY1PoQrLOkK2CJb+MVBc0wWm4H1eu5jI+pzu/KU1Mtdkn7g9v6Tz1DdjJhrs
R/Ol0RzmBVNevNB9FuPMRBNdsQuS4KPYpwJQsr/kek1/M8nZkdl8KyW1gvRZE0vx
8mHMQvZJy1fVnqNi/kd+cyZNZRKkVhFcdgh/UT4Dc0hLJkzqWrXXuipY6c9+/gmg
LZCIlggXxBQEn/4YNrrqtMAuIxNWnvhMWxBbRLSUGlRzKg+jiq/QaMkodb2ZohX+
iLWlAPiIoPbSTBbNVFzxpXSRX7rvAbRwnNSV2HfdGh/B9SW/auMsEo6H+UtZfqgD
odh50POHd/Dg2F+m2H1ufgNX3agv5Z88s/gjUxtOmUoZS0L2rLwDKQYz0QyQxg/e
5X9vrvfc4ksVzB1Pz6DqrB2VQ58MKVSz48L5g2onlDI100s7DKIWJHAx8sjAAJ4K
AjRIKfXwi62bfRbJnGkMj6YXzfdtHJO3FIVkoZIO6izDGq8FE2TX3qsPlf0Gsks/
okFi+VInpIWgrB0OZUx8LkhCPvuh/scGM9kQKdZhjLqE87nfMsozXoGH091fg2jC
cXiRM50D6yHX9EDs854b6uouyen/0/XvIK8/vGFpNb2a4+md/M/LY5sF3QcYzM/0
c4s3o1eSR/eulbD2n97Srsqyf8LT9K5Wegoi7+YJrwY=
`protect END_PROTECTED
