`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xil1/uG0RR17zlFWdF0/ZH3V4/y+iXcP6gLH2qIAIsf
UNjtQjeDrkKtE93GOTF7T2zd4rFpnqVDZJt+XgHMc3CQhX5SdwwXgpwx0IZBuqzw
tpgHziPBTkvpwvrqrTVN7qeZPTEOykoNwIVg6vMri2RPeK6GNMYBuVhFFQyJe5tz
Kxs58GktWDSmsmuxE7//P9ruThzLankjzxzIm1YoVpOoJ4JSr4o4iDHVXr0zq1c7
OjUZHTISMa4fHZAIggN0TyfDTeqtT/eTUXco3H1CtLmlQ7J62X6e6fYUeVcIkhHP
cR0fUs6XCrWr5h3FP0oHMg==
`protect END_PROTECTED
