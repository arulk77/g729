`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rPfN+/7oEaa3Gn/2Bu/2iXokEGBRlkCaTZaGsJaAM4yeMceRyhHJIGhtRjSrQVle
yxe+d3CcL2cs0xoIcOWfRmmvRCS8Oge90g8a8ydcZL9D60LVzYjF+RnlmE4jqS05
iTz7r4mZOdNVuhJTHg0JU6TK/7k3/Zx8qs3mMk76G1gIqmWXjusjj6LTouVYFbbM
ZHCnUw5IRSQHPcfJtTCATH1OjQJwZoCSJkqs0pwXo89Z7OCJjlFBURDr8vK74LJN
NzfqDuKNwB8Al3Fu6sEYZKJL9FpOnBRgaTV/jtPK8f3zd5xPMBlAv3OdKPSx1goO
UnZnGltFsKRYv1vjz3zpghTEcXO5twGRZPtUftoIG1tLmusMBZfJBeEGWFCk9sT5
Hx20O2DyeM/p1h9baR2Ai5ufTxVB943VWegojFFZYFQ=
`protect END_PROTECTED
