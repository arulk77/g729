`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
S4Yr9XGEx4jbNmrPEN0wKDf38aq4+2N5qBzssEEPzcdjBckGk+Vrky0og/dTxeGQ
RdMiANXO5HdOa2dQma4RH1yYf254/3k6K1EHttsMqLsSQ5Rg6zqCF3ItK92a/tss
MUrq5r231pw3JSMa0aFyv2zCPaXvSfCzr/fYxXtOUK+RQ5sbMGvu3ACS4KHNAx+S
y3FuhxSOSBFyDe0EpIXnqxWUWzixZGaXqm84y4V0Mfllh7NQEFAlsZyn8pI3xEAw
CvOU44TFxXEoW83aLPTc3OFYsgeXEpWnh93SOWYsfJ4ZlN8tF2naVtiQOIVlYmln
kXHZigBjJLnFto2kNh/UrqaSHYCNslq8Zz3TbDDu4TgFd/QdVIzKgOgscwI42GrR
7JqUbb+mSJmjR+hwTUcGng0oDj29btCul4waexf70boDs0bf71IgYY5T0DQB32Yq
Nnc8od3EbIcsGiG3mKasiOt+hvX6Sf7XxibVzaYA2FEi7ax7i5oMw2dwimAvQT3d
IaZrs1KT00n/ENEanSEe7bwXb+H/zUS43LZCdynkhyFgMvyhtGfY82jIbV6z/lbJ
AYjyvB9ja1gEQMjTNRjZDk/h1H0X3iaGaRhW4qn5ljQqFAnltpKXHNhdB9b2qjoi
2IZcdUZjSYIZGRTKjlkEZ7emWDOwmj5aGDLzglduWGzmJ6Pe9JIUXW+fuxZI4WS8
/YLpFNnDEgrJaUd2NeedLi6ChIGsQ515S5LDF6r2Dl5vqfzDtgf62RSDfWVKviTQ
gG98bQ5kvVfCJl8Bjxs1XrKRVEOtG+uvZXKlm2eWeqzINHDhy49xNuVGTktuOCYX
`protect END_PROTECTED
