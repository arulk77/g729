`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
U5TIwKJFi919jRNElPB9bYDvrt3D1bzzbMWjZSvCbn7e2EFjHlP/ciQ1uoyMq0U5
LCO2mB/xtzIF4apHBwWCGvh8omtEoP/wvMkWFPnE4Uf/vzu2iXoGXk7GCGxcH5Dn
P6HGHqgDXjneHjI9WgTkhylIgDij5RoZdAEZlkmiRN9YVLBU5s0cwZpS3LMUcA2c
L3AZHAex5OyhUUVVyhwjTy3+KT4tuSjd0VMIrDiuXLocpIbTdjhfwXivcPw/46bV
oDUTGY+JBfQYxXDPq8EKkp88PkIKazz7yzrvC9EYZAbPk63vh/yvcHjVhmI/vs6L
IyWXJ8OgllBqfSiZc4/mDUOWPAdpbP/YBqKJPpLIB2qXJ0Rce4xU6BNdmEB9rOKN
Pz6Sv2c4EtsjI6XszqoEds04mKVOoItkbN5r00fCnj4wsH8fi1fI6+TuxDpKQNx8
966JBcjsAs+Fjxb/o3uYSQ==
`protect END_PROTECTED
