`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNpDvMj/nIo4LOe7/4ulSS0hkbUSEggOJTADSAMM1LVN
TTMIVPdR7uIemASljle1RBJapYPLvXF006v15+WAle53o7Kuxp3lw68aF45jh4Vw
C2aVQtC+BuoDBPwzXJYgl7cWYVXQwJe9vwpoK5E+WpfId7pqYx7ZRUiogUQXpOXA
SpGWBirBiLrwfJ7GPlaIzm3UKRmF2PjKx+tkrwCigueCzSR6x7LH+NfDTDqQ9RAZ
`protect END_PROTECTED
