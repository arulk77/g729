`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+hewB9LAja0xTYohsFiYjhhcMa5Qm9tnHEaYn21WngMxJ8+ZFWCu842rQaK1RxIx
FD2eWYS0YrEiKt/1d3yvMBOk8vLd75xeyEuK0zoFuc7AQGMPCX/2ZBEEE79H0bDf
A8r3aX7RfAGtuCTnfHP0fZz6L9qjaErq8v+TfIqUQTKHECr7h/9B+sGi+EjBCaTC
rNxTHc+KQxfGPU0PCBHs/0nHY8U5hbm8C1cqpsPehMfBuApNZUu1ayKozSoyawyM
L5XkTs5E1jXMiPT3kXRqAVjGv+jEEfz+0gmqzWzOKHfKHMMVDxY7Ue90t+C7xkTI
HxjUoNmobLL8gujiwmRlVcCSNhqP3KMBkI8ylO0TJJEjgH/xn6owhxotZ61M7JXe
z6EWmcFG+Qvrjhou+e5bqp0wg9+7dIq0dw1k+Ei2c/i45zCoYfrOrphy1Oxv4KD/
PbWNZ1hea3hxmFShgJZ2XgcJienKq3T/yJEC3X6NgLlX1E1AeRcgnohCugYsy5N6
q/968o0IPwQ6SHmaXxUxQplPJ1nUUER/+QoUo2fETnytHMVN1+0Lg23jxWjaEbwV
b5vIN0EDbFrQmFt/ntPuXA==
`protect END_PROTECTED
