`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Bmt2gG/yp38OVZu9soSss22al+0B/hMHCHMVVF+zMy+7STRgktUXeSBC8YDkpb/A
PmBLHs9o9Yigdx8/aY8TSBZvQfCJltFP+okxJo+nLyr4QwoH8WqMQpVdEZF5a/nF
slJxC0dz6Cn9app+i16QDJSa/aEGUiAdeZbXiO7KzE6sN6Bc52vsC9Dw1ENHnVPL
`protect END_PROTECTED
