`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDcZGvMYfNbnX0ucjmhj4j4+frbfYEUUt6/m2+4lAnzK
UHIGllRZmUiPQhj6KQjKS09c8azul7UzfNviXnAlXlZY/8RthpFHTWXM0/i5lGfD
e6RsRtOZwnh/BdZsH+sL0bt8EbYlVJ8d3Oq2QWh1V7RMXKu5HYf476Si2Jrq0Xye
6tQY11LXMsMITmToKuIv6JsgZOWYh/u3ZDfYXtuFEZlLB9s0KUH7ds8KdRrD/zp7
U9P29dwXof4K7NG5zlzpg/5b5YhBjxA8p/jD7VJV0uhtX4AutdQs+nhy8SP9D5K8
pVVGgPalP8RepLlhbba9mWJhx70nx9vTs5J902WMNlWE8+VcTk1ijleweeLMVNN3
cLzXXp3lLi9Etp7ZpiLkgaiegFN0jomnG/kA+ZQt8FKxBnzlvZgGoNVOrZ6Azk45
T0IMHBy48QiP9jMFywxNemGnyKlqTuwYfaQUQvzpBUKzaTSmOvA8AwMsAxVS3vW0
17oSRMd2HNVt1zPdiW++qqsxcygHPgMHl/ZX5u6YpPEmqmHGPeuDVzDtpw7/Yqyi
KmFhQB6p5qcI/lwBctyCiQ==
`protect END_PROTECTED
