`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK3V7zffbhvMCwL01t8QAw6yNgAXkUE92ivfmkW01F6s
dSqkp8lmP4esQZfOc84ZKPGyaCCItqavfMuyggWjdR40ZFEwAcKuxMrJ4Wlm9Udu
pjo6u7Ay8YKdULDeKF+AeUPPfRYDm8GzNgxjz24kFMBYUQZMfU+2M3oCPEajvvit
+qsYVzH8Z4/DlunEnq8vyChyGDzi9JpIHE0E4ooiWz4qTruUiTSHYI1eqdEcjqar
`protect END_PROTECTED
