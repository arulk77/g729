`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46mZvibG1ksTClHzzE/ksHlHphBOgSm/Z5t5myrVxZ6k
KwGE5DNVheA2M8eq6Hea48hiGV8V6tLXWdXN7+MQ3MdR9KKfle4pgQOHoNE01BdF
6kdnfyLn530SH+SlCu9Olcf9OzbkHf0NtsUNVxoG+cop/ZMCOP+U12WI1nPyZ2Ee
uknpfEVGobyJBLxRp7bPa1GO10FYBQ3H15wqCEVzrh9vRe6b54CmTvO+B0DrKQIn
Eb14rDSi6oN6PYUew9qH9IiI4MrzE4MWHTl8Jwa/c+E5+oQZu3FcvT/jDJZHG2Ce
3VGNIJdz5etEi9C6Jea4qKWB5DbAc+WsfBIxpTTEGraMcEmbFrs/9MOz/uVpeUb9
hnt//L4AKQxW7+oQzwokcA==
`protect END_PROTECTED
