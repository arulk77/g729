`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNdUKXkcTJicwsTn9dv0UOD7zd0U2zGhzLWB4/9OXvD0
C8Gdi8CsNENjYUZCteRRoRQgUJO6+eZ6nPTUWj2zPIOT8U5Jyq2PGxRaR4lu47hy
0l/xefL5Wly02KAdCobS+04xv+W1ezL7VVsFRJc3aPZ4lv0iie2Sa9Y/Joy01yJb
NoX5zlOsHF0mNaZsurVJfIbZyGthZiVKi6DFZe229S0pREu/8E6aGlMMhiKG6cQy
aRUt70w0r8ojsSj/I/FMJzbsrHmP877+2negRGSS2eN6hmjYvWwH911WkzK1fats
VY+ygqQeQbQLiDmtD7G0UMVV3QIdnJjEsTjT/BKxZWfd6Vu5mVVqW2SxiWoSI5cc
VNNIgYIL8KK4iHIR9OKnESFh3V5JrD/smeOKy7uMI8pUPgKZSpyftTj7kDKBM9UO
UOXPl6vPY8RKJkm4E9GnQeMalKmyxKVKn2HuW+ju52tyivhOL8nGEsI8Kd7HS+g1
hsRqZrQd4XI+KhzybbpZvLH1YmuBmzQhsbLYtHbj0ZYlSlrLmbZ0kWVcucxvePpW
79fva5pmHWJkctgZ1sziJB/JdAB4Df34a4G+COnc2D/4CFfjmX8L7lVPlfDx8bIS
8zV35LVQgMqKr13zNk6LYWv6NDOnuyZnlr5DKz6Yy2tNb8OJQHNaWrFx76kg7o6c
rmpUWHaZJiiU/A0QrrL3L6fdhsNc/3xtgW3js3CqaZamVfPWNSm/g3tQ87qirhxd
9psKlVPy6v3TI6TLvmp9SsJmVsJGpYoIh26UiE9rq6JxRyCWVdUsW5G11H2bXJ0u
vWg/Y2K1PrWzGFB5DXQM8MrDkE0wLM03EGL/pozxPI1UNcyk6La8WH3I+GMG3zwm
Vxfj6JDslJAyB57a6DIl6YMPOaef0BOflRsxBf5qm+FU/UyptjUXmjyza8fEtOjH
9p7rlLSh9n8/i6RQ2lYKocmCmPfhy5SPuNi9YA/BDF2+fogU3xOXuv+YwbNoNJnI
GKkm4q0hEyQicX1Z8Scj25eHvCtcbh9ePInXpfQ+HftodQWKMn/E1Mwg0qiUzUYR
3vjTxe2/kET0ovaK1rtdtzx5s2E1jvO+FqcBFXk19CVVJqunbbG5ACuzxinWCwDK
IGiUAqGlbmaQ2TsGSk0fLVNVI0M7S1War2Ygu9lZ20w4xVqxEwM4vqbdRkSTjTVA
cBPitCNj6dpAgVar0MuXaSKhjbGV5HVl4jyDBLSbSeYvu8XiPA8Jfb49umVxV3KO
gJrGuCWWO4cc2mG43HymRKjyKciURZabBt/z3cDbQU5xGg4d88qRuuYXtSf/g8Jm
IHy35L+nYXNgSL1cxPyUYg==
`protect END_PROTECTED
