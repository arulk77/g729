`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCAlW3J4h7FYKLsPaLPS7zEUryaIWjeT7v2WYPufqpC8
K9WGWNP6FYRQRp92Z7lay1X9BfeJhtopM28+5/xueKdsrLjESr6VIETPv7r446qI
n/Nw2nPCPOIPTLPw9hlLGij+t5E/LgUmxHsx4AjVrlGUtjvYRsZc1g5fvVXdgkF4
2R/NDEc7nYDOxY1CB9WD/wnj0Rrnh6VETQ1YzKsSXSt/oZ/C4588tnWSkg9DFNPk
5bA9DleXb/Xbp2E01swf9cYwEDa6gKGCnQTttX/iPI35gauu3XC01pdkdRT8amwz
auB7iYn2ZEtWaGNWOqbyS8rgShDk38Nvn1VEDK6+ckdlSvTs7ECLyJhuHA3M62ZO
GCtJX99fagFq5vLnKV/Jps41fBPuo2yK4nfixmqSIbylBlTLiq4Rdq6hASPScfbo
VFc1qoOvoU+98YBceAhoPCTzC6+kqSX4nOeb4t+aGIFwEenxXTliFacPT7zedEMp
R5gIm2SJoFLITM8FwZ/FITwyiKGj/gBc4SYPUOz0WKTxcyqRvGFNfmzwCiPnTfy3
qMfWnH0HrqyCt4piWsTLYPFeP3YHHUTbsj1A8iv4TacSIA5Oh5g3tkCxJ1lw+l3I
zk9qRpPYZ5O9Pg1N1E2bsBg5mKl6mplx7X7YzDzipVfeZMxT72GDa9Z+QUk/XWhJ
F3mYz2+K3OmkyyQM7NrWEEsP5jekhJAo4zKIEaAfBCbODkiT0sHzhCbkPLxsQsl3
++l5jHpvIYJjnT4MkCK1XaxyfR+KgjO3ifGHj7WPWAvJK3iVthU1/UcK2FXV9idt
qYkiRozk0RiTS1CQ6lyNX+RVHJEkws3FnqLQV1J/BdcXIN9wLbjmqPxap8MjxFUK
5YZa/k8dgxqkyC3wQQ+/91URIl0v8mLmtorAr8Iog6lcvbMQIHSCzUxtDmcHsSju
AWhGrrmDgl9FFzXP0lXNn3xWNqRSgeiLY8R/mI6fquSyaZP9omR89Vp44unKkzNO
qHu67Xo6YYCcz6m1fg3aBOI9kKhzv6fZLU4/QODQcdJUmAFO5TeUyGfreGUpDlnt
Nqtq2u4pJDsfzrlzMKpx3LIsAqiMH4DmmD1H54PrCRRbSA3nxDrds6oPKzY/YnU3
K13rilwNsoF6ZHIiAQmucA==
`protect END_PROTECTED
