`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9PMRcKt5l6bV7o0RiD3qVIomr2HfZOeXY3qKJILVsNkpEwbVsYPAQa7TKWsTy4Lh
9FtLT+rMBhiL+GYvkvD8QGf9WV2lWN/lMUDgyK//YXzbRRJn5i63378wDgG83pVp
VsDnq9FCrCjuEEwfUqah/7i+JG10Q92Uz+VYsCG1Dk0E9RFc2JQyCN24VvbrCZrC
eQoy+7PnWqwGosJ+Zk7cmvpz/mp5p5Ygsc5vOGYHXYEy6eaf1D2Krt+fCplw1udb
ON+IPKO+dt414c0Qkbb/alzaErKTPUUAV/ZKCxORI00=
`protect END_PROTECTED
