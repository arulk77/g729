`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C7UiMzvBT0J07KErcpGAuPAhtEXb6FKJMc0YOhxxUYkP
cy0xbsQ1I27dX0zzfVlmPOP2o2A9hL3QArM4STF+NUPThRlzZNmsxaY/3bepIupr
LppY5LX0JV/BpzmYwJxG1KHexJTKvsDfy04R1Zj5v2Cvy85Ass1gcIYOx0zbF6gX
QndiidpMbtUjI24brvhytPvyL/IcrEN7RpU3gzmim8Lqr/sOVVq9cqr6a1rWmOEP
yRmGTpM7G0L470c5bLqlUP94feLo/9Ch/iAd8XDtj6uYf45nKh6XDj9DRLPJVN3Y
r6t/2LISkqpF46QJ8xwcC6n0Yh6ln6M9smOSDE7xv+IMUL2OjZ0dOVE6yjWvEDiO
+rm+GR+OPGBmOiCsy05vBVkrQBxD5zQsz7topGGydIOJSe52ufRgdTuqJGYWX6w9
uIPupziWxWhJGnlkMNO2aCMFeU872bhtNtXwTCQR3ZIKlWGxVzSRzoF/53HgN+XO
TPKeSv2lQ3ve23C2OjcP0W7MwlwXzS+B/SErQ4jX7RspPPC76BnLPbl25iQxnVgy
sPBJCUsnVvNfeIEOXGVaF79mIfLuQ+Zi0AxbE5Ubg5hoHkk/xCFyT65oB62+Kpq9
NVqSAlT991bzv6/7fEmYUhWaypYgOwu0xw8QPNKme77jPeUuLGcBbRcQGvXNIze4
SPBFGYD04xkVTPewK/EHlQ==
`protect END_PROTECTED
