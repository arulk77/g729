`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLKk51LF2pjomnjfm2iL4s26i1JP3cz49VcFgXC+KFnd
rNx5Kc7WKGxPRnre4Ovl2LRLEz4+I9Kdci4cbpBZxaC0BY8Gst1N2Ir5k4OT6Gzr
sk1Zrv5507DZoP6hXcwcejbiZ+QQa/PpqVWfw1ZCepcIlfd0KL2GVxWoEQ8LLDBR
L5jOcLDbAEB9iSkXHLDwb/OyIpcjZIIuOi83fl35YWdSTBoMeSozAHJJwqaawWjt
fzkWNHiu9GVzoZ2fmdzh0D3NFXe0LGCsuLyXLIPHJE5L8RkKrA+ypJIHVY4IDizC
2Slb7dmcereo5pjgaD8K89bkn9H5GGAn5nFsX0Trarvzl1rsC8qmPijWnsn5IxPh
3xJk0r/qHL88d7Xj0Gz97lheJdI0XuNO6aoL7naRpgBHrUOxM9K8pS9Z8MVIJ7XB
Enhd3lPyMCQf74A7FpTS3bZ3oFPTTbRvrl0VobqjEjMl1VOblElLdl7DkVjNIiNr
sTTsaZStXe6N05qayI7Zaa0kU/Ut5Ltyl2jNFE3E1zl9ICrs2/bifOt5iyCx3S3N
yk3QOzpeOk1zNMvtPeR9bDABa+mAVmaLFIKaaEBBJdg=
`protect END_PROTECTED
