`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu411GXFXf10S19qonzLeIJ+a6lNppPUMLpj3xKECZfMGt
ekMs6Xs8GhJNRTbZJI0X4mAB0rkwVWKWjFjWTB6N1uo/iMSxI5nOsOZE46pR7RxO
RSc/Zl9v0QHSxBMrVsOfwkaot+01eGEs4G/BfGTNFblZJx52y759orR7RvGitPWL
zFSMonAJecHCLZNxO0IUEkV1nk4/T5ZYL9g0J+ozdkAf0PSdmB5aqT6fWFfxXOXA
JT1i5P+2sGrHstWefJSkltRD8FxM4dI6w06kg64VxIeaywkhk8LRtatIztkhxMLF
e0aulpCbox0Uy6XpLQ81aXThXdvJlCtyGOggFeFFV2pqPPLywkmSXCZc04HIT6++
l7P9n1MJpzIBkT5NuQouVA==
`protect END_PROTECTED
