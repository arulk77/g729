`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/TruWx/JGAEOQle9H/xhnOMc3s09GYTmHzqrDh2bvZK
StRqXfZ9OwqXDwT8KemFqpc+Rn4r/aAcghbiszE/RY+rxLp/xnwbPVRiiQmKk4YI
Zei1s+UZ5zVhiG1yF1U16UfYe4hgzAjpyuC7gJRuiXC8BbnLaaFkK1a8fcTvatGH
QH075P12yvelk5qe38Bw6ziouaM5xhpFcUvAfGUGDbrMPhmQLKtZigcHse0qS1Vl
pNPD5Wspai8ZwzOwC08cxQ==
`protect END_PROTECTED
