`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM2oy3NOWK5GrSGFyFML9gTmXKW6UtrircyF4fFpQ24B
BSkJGBPdzFXPpWOi5E6QE287iitnymljMB7T/LPV4EZGHNE8I7c8Q2YZkiXtEmVe
LsaerGwMenBYcOwJf+V2jeXFXQB8ddWoiqOOSjt9z6sEQIYu4gciFs9yHocYQFT2
PUaTXfwoKUVexEYJUzRCkHbEPRNU2s3e5pe1ciqxOgNMub1VSM3P9ZXV9pQfdlIj
7jV41eLLptE0nXPIxgKlR4O9odVdo+V7RNFYzeSIYuw5UtDAYNvt5aOqKQuQ8KYt
wHAnyfhJR5c7Z3r79mVUG1ZKwoPbXo9Mm7ZaVHAStAsU5CqMU1bfYVc5vwdTmGUV
1OpH9kGbSeg+XFZ6x2codpGhsI+zFXCgOTUQgVHovXQ2/FaEQefFMgVi7aMrhitE
kvGqF/NoVr2swLwJDYpwCXsLbdbacKbIiSzIwRYOe0RZqeARuXJDPTGETwp8NZ5R
NHdLYHgVpFa0vqKH0S99T/ZMEEKGi80nBm6k/Ck629PAtoHgwnceSKUrbuxfiUrn
`protect END_PROTECTED
