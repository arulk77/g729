`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43/xHzkNfmT7f2iVUxB6wzzkZTo6kaVUO/v4LqnX4qci
sR7rlXLpLg/8/2Jc1vx03GMKe90gaAiVqeCgDrtPfV5RPbfq7PBHsBIaCHFwAy8I
wwIdiCRgz/sY6JL/usLIkdRKgRnlX/ps3rkS2DdTsHQTHl8A0Yw+F3AQiZK3Kgmw
xvE/LsNtlC0R+oZhIZNI5/x8purcXz6fnrL+scRA1tNVPp+NbS2DgNsW+qOEIzDw
u7g+0yRtukZb22ehALwYYLME1NDYaLdnR1Dj7flcus9ywkUqtmBoz0VK6uxAG2Fb
TyJGBCnCZrXvgMKINL9/C+WlSJEhcvhZX0mM4L/7ftlVxyw4Fyb3oytVTq4+Yn/q
/LcsIeDMGYPITKEN/2+23g==
`protect END_PROTECTED
