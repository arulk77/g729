`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RGQQpsB9qU5MBDVn3OzP/NzbMW9CutZMGcTyz2Id0zMpAQpSo6Jpyt4JB4UC5e+P
UOFsbADAIS0elUr8aOC3WhZ8YOFDrHRpNrB2wCfYGee9HPrStw2c4JyvcbPnD+bh
Ko7/Og9O2Rt3c/kH5BrN4eVP2pCS8BhCNADkOGpQKv88FPZl2wUpDaMF6chQwnjx
tiJQgi8M+gZC8sZtNvqpFq8708FOdXW3SteTSi+nYyrwi/qy1SLwEXt4ovAWBL8L
D8c0Y1SBTxtp6GShRn0PhUqgrMu3KC3sijmC8kP5zrxFhZ8rKZ9UhTJRYufNYOCF
`protect END_PROTECTED
