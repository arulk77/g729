`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RXnyE7veacffTNfN2R7SRchiUvkfrfyqv6xjgO1jdGWgloMcZLjkZP9EMnXiOrJP
TC1HQnO6CqFX7hfmjZYP5Sn65gKlwU5NXk1yA/ys9QfffJJRYDaynvKapdXStIja
9yLqkvelKJEezRXq+buEFpXt0/jzkLanaMYuzQKxHlIm7sF3tHyGfoUcdeN4Zw9s
nhAhYP3J7JAVsNGE7jqXl0o0Cvm5p45J4pUN5Rf7xuSoo35LEJOZirVynoQWwuuQ
aoVAfUpQ+gMndhJ6IVjyoYRND1sPD0/se4c7zZAxksWvYNtqoxYQTAgUyV9Jv0Ah
/WXyPwQK9g2AnK3OTQdIGLMR+2MHcobCxbVOGePFIw+N46CnCZcG811dYTUQxUpE
UeQd6NDg7Pq2fMk03rm6VTyoDFuPW/dZQTD1mmBpKlqM5hh7eSslbPuJgqOCY8NC
zIl/Tur0SKp5TPi+vIr6RuzKwhxU4qruaAgSBnYG1V0=
`protect END_PROTECTED
