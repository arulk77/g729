`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLVAoHf3iczE3dKT1wNm4x8VcnYY6JUPv0TnxPajmv/p
WJS8NZXclsOT1w92bsIqbw2eu/aXJPLGp6aLCOZwodOwJOCDE6UpkLEA4PwZEl3v
mGUp2UWmD41BeT4dB/iliUcACcOnd9PZ6BSY54I8CymGl5LB/peSahBzGiDRmnJH
WQRYAKLulZ1m1Tto4QdPWIB8oKFTLj4gYh6uB8OJxh44XYJoUI/jmNxWgJoH4rPd
baFPrA+1IChLaAHMrnyq/s5+yykQbC1mgOp8r3/CRpaliaWdyrOWLkbdR35m75Sc
h0jq2wYbIHdaYxpq1RTm//h6uMyX4XaknzMD9kNkGqoMT1DqFj9Q4DAQ55hSnjtW
aMQGCxN6C2Odj+2uTexEyTGew3JsI1Jv7Cd21Dmtdc81RFjxphdKgoxBXz99ohQ1
UVqkQCQ4lRa6mJIBgXfg8t/6+YXhanhDk9FytyuDu2qmU0ZlE03ZqXF7MM5YriGA
mBboLwkVKvms0qS3lg6BTeZuFWEWR6s3+RGPlkOqJ7dT3+0yHWaQNx1sGFzqwlNw
XNi3lvKXTtGjDLzo8zK4hk21QWT8vpJ2qFw1sTXZR1drOwDLRCHW4l+Jlwp3LkFM
NQKdQQYC1sfBBa9YVBIa++fysCgy9lIQyxgA97J+1GVs89QbmavEiYGhgi73gWi8
d35nZ+IUJYiTOQZ5/DXcHgZCo4uWb7F8kQC93nnlHzZlyS/4UGjzKD6XmUrv6/Ej
KfBFTdtXPAY7nn7g8oa8Zn9dBtARjgDn5x/UNo7iZ55dDyei/TbIOAh/G8Vd9J+y
U6i6v6QDlt0oWhdrTKqWuzKIFyH5uF4NXA1N9GNidKY=
`protect END_PROTECTED
