`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ0OmqQ13begv2W2MSyC5qHr+g68GM2C4NLNzZjGxYhE
YyqMCN2ajWNYjmFC6zClh0NfupZfB1Q3noQ8FRODCYHTFFGuGlDDtWszKFlw7uVr
EVtgwHfua7i7wRhbZoENDfC30kr5LoTuIwLKoftANOD5wf/Dg/PZqogQvAVxggk6
se3VSIjlDDPBB5H9SeomSpYOD6ylvEcgeIcIh2KKgt9RBVbHdsJgsmXNEeocXYZ+
xsQ4zOrBHjGHvnbbtxT5Bw==
`protect END_PROTECTED
