`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3sELc/lpwlgcoWj40fvp/bbCE1ITcDgnVD7d1AfNyGnnK0KJE4rkqr7JCTHQXK1i
3zDSthvYmJr66CQi0EnljtxvQa6XSQq/Bm5ycE4iM+RwwgZkyY9WsJnUHTsaur/h
llqMh6+aTDFeRaiFwsK7PovF7TS0flgfuZS/dTFCqXtC3/NTKmZLg5R5ImI1cQEq
7G46dA2wyiJ7p2pmZOxd9SuSqohU4Vrcz7S6Uzmm6N4wPiZGTAAecJg8oEOeaF5w
plH8umhLu8md7HL11XzqvZ9S9riFMu7HXQBo2o9Xy7Jj+Te1zcSgeBgXd9RyyDJe
JPmMQW8avFvJtg7yspKoteIGFRguKuCyp0nxy08abZqZEcja3km6pbvKXcyeGVux
92YJxAUOdnyzGDvQGH8DKltoH8D7GEf4yXGlI62bkRATIhLuoald5vE3Ji8/CG83
ITQSUY6greEAZhBX+NF0KvodhHDs/UwnMwy1SMCddi4hJWO4M1g/o3Uaa8AT0pZP
HV9DzuAvIpvxcaYvojrqyHayVOoZqBe+/LCyH8GwyX6BjyX2dkyMvXjFQcQ1wt2s
jibVBHx3nUmb15Ylq4iU5oHhBt6uJBse/LVx7NZwsrUfN+dxkqqjnkD0+Cf927Ds
ACiCqyw8+uul7lNjKeywUe00Be8R1xcg5cEjK458Qqzx4aOUxRKIbgobwHD3WdVF
RG211RQrpF9suQQ60PFqitJCv1YAiNCAh+Ss20pY/WMJgr7edHkfEkgwMbiCNVzg
Up+6LIu4gB7F2W+6ONc4UTs+mkidXIe44nmWCSkohOVJYNRFF7OtGSMz8fP2p20X
7T4n+e4flm6zrRPWRHWRzMOmwCfERsh7diFU9zqhRKoBVltuqcWWIUDXI+zisS5z
DSAy4W9Q+Gc7Ggurmpm3R34aoS/uyYGe+XEA/nh2spzmYbs0+u5EqjVLUgVFQUDS
RJUasEBBq4AbxyuKFpcGWlAhLNP9U5/ZAw1kKxsDfvspPAG0ADmKA/wB0UIlo/Ak
fXZGZgvajSB7CPVDiPj1Zf0su63ZeJTyGp2Rin4At3TNbHk3Ur/tTmTk1uhLp4hy
E1z2WrCpNpbHuSsj3xzmR2Z9hyZ9c2QVAUkxeYAyF0DSpZUHkw60CZQz/FRIL87p
4fX3D9aN5whpu1nvj2JYN3t4rv5gm29UlDjXMWqdhK+M0kbg5xceNvLz2k5VYJ5o
Nhvew5NOs5t3yN27MtjoSDfVuTiAjXqrXSTTYchuGNd/44YWJ390XBwvtCAVtRTG
UPo2fHq/cubauNOoxL6R58q2DBzQ7whkxG2OdzVUWXu6qMe+C60XkbWZlU11uzsc
tmcIrSWq7DSB+bj9ob3ym908Dcim031cZnBV4re3xRxTY3UP+GkG0Djt0SEJZ+NN
Lp4cWuDmCLtcbQKT61i4HBmR2IBuJWgblG4JDo9HkTQbcy/7RhLENKBaBOEkSrwb
i9LHJDdTXox1v4l3Moa2MixJrLVBfFI4r4qSWLpjTA+aqzd0swm21khOMmQNmbT0
W4kntasSjhM5kPLZzo71kkMmNBUd7WPhBi12uWJVujlnHctlPU8JQ72sFhZDGgAo
aWhjEbj/68PkyfUW7DeOP6AGw/q4LVBAV1HZYIOVpLbKBjEiZRRJfZbBqc+oD/Uv
2X/ssCxcw2wvlGnLJ5asS+jBrAxCNcg5SiNZDvuJlbDuXu/c1jZIl4CGSdYeDGfV
Z4Vv88uNI9GZtaT9BSl9xJzFrfcyPEZb40ugPQenCLad2Wv+oGP0+YZbSJ69Ulx8
uVo3hRUHPJ0MWnNH7uvMWWn18gqCZ4KfJDf+FyH9VeWeUv20Ptpk7FLWcrH3zryH
x2+LMPO2QRyVcWQWlZkoGYSjw6sLVdRmpvpSkUKKU14Zg2wT8PyV1rpM8+huwTj1
ofj10C0pQQxy3U/Df9a5oYuDPrNt2kiE6sguUveZBlUZLzNTsU+TfcpAjOLM+Vih
H/fqI0+G0HrVYCXMZG97RVogvPoerUA8wKp+mNYziCMgoA8dxfajzvT380dwo1DF
jYJ66QHUzyruizlaWFyg2t0nKdz0RBecmekcr9a2oC4T1WnjeZKUBlOWYFPepP1H
oigLN6w2KLlF6pIrWDG6JhfOzUch6qIkaZvBZt2Yp59aQg/8DwrAB/hJo8RElX3Y
fA55ZwKPMYSE7E/4ZKUffpgpXRU1jIz63BurN5tXNIW8WiN2vx/I2hOJbsJsq5lM
jmK7A4YULHZU1X9c6mvyZvR0q7VueUsqGXS37vCojiFJLxH2gTl89xMwosGx4s8d
DQ2c53BWVPom1lKxQyHcgFEIuPHmnQiEXYtXYwBgYaZ8xzeDrGCghMdi9hZPr6wI
0eZUBaF6/wTiTGux02+r+5/oXodc3CvqC4CNEMKJLosXDGxbvoCnxaSHin0Kk1/a
iY+HLO7eqh/9x+RDAJBHi2xvJk6c/yd9evR3GANFSdC9v06Rws650JDPTPF8h2PE
+AYCKCrqZFaf+oJxFWXHxz7Orr9+4ZffdB5B+tam4D0LA0pR/pEwpGNIdym7QeRF
MttX13AQedcY6IIxY0D8nCkul69BvqMcSWa48Suq97MFP64PzsH07UvGxcnMVagC
`protect END_PROTECTED
