`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF+fKz8ZDUDhpYiAvQc7PteDGWN0OHAWx3A/SC2WNaK+
zX4PM6qOFoVpaJwUCndwkWa37m/IXw/xuzS/f2e7xFZPLb+fPVT8BB8K4PEymdrL
XSl7xgoYmBTndNCr7NSGxlAL2pAsCBX4BBHPdSDatP8XTA899MLAywaGlxITaA2d
Y6PcjnxL76xXX4kHztlWoKX/KuynrdsRj4zjg792VuhSkoygI/Pzp+99054+VAzK
56YoTNkb1w1PhqaMXce708FpAzBMvOeLl8I+PDufqc8swYEbsVV5ImIL6iQPkJ0p
7JB4Te+ev9ZvEdNlK6lQoZwwd0/1l+ABpFjGRoTAyh76kuKKt5+x3cKnX2Te+YK5
fsJqwaBFzMioqAI7RH85FPVLa4htZc30MGKX7QmHBk+GyPPsqEU7leRqZ3MNd2Ir
EbTPRaY38+CT0xRssTJ+1paOHW5NapWeU0aOUkvf4NkwnUVs4p2xuusKZIUbW2a/
dwzt8MPkodng+YQYCQH1imkbO4RDi1h9PL9S7bHO02INTHvPdjwYM3rtP8HXTd7S
DqZw+PUc8fSL67kXTVHPAQhAu0VhRCeD8ecRbFAII71G0/feTTljTGs/AbyJg+gy
G8/9th/JlL9Vk4d4bUmc7Xes3JZtRFDBXWbs+oCZFdUYdqKUEz7MiMhc94lp5qCx
Ek0bDuAxTOBOi/tSOmSiJrFX2iztaHufz7IRfUeKyy0Qm38eQT6Z4dODPlAgOiPL
MeI+jEXTdCJqjzYswumZ4TvXe/u7i+hb9psn8iWhrqUk0zxt3Y/5kl+NXp3H9dFh
`protect END_PROTECTED
