`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAQbXxgZtCyL+BeO55x/CBoMNRJAe1izVYHqlkIttVbrf
uGcKHmHo0730BEybKLGLVPP89aAQNYNDShtM3SkB3mwZv0Rac06svNEQyztukUli
EwzEUEkCPYyUrfeJeNKQQjM27isfb1ekngDAHJl9mRBrJCyYtCDsCw3DJ1UGeLSb
CG1EY0rGlgjWFE9c0FQ1x74S7k2uk0J3md/USbMer3hyyd6fn233XoFfyF6rp7pS
zTVVFcxIFbfKjAceCeeYG5Keqmg5k398gFdL6PlYgE7eY1usy1ciQN6tcfemIvx4
m4fiZN+SuUFqzUbtT2D71J16EqlQ5RtB+ZpfHYHgXjXruMheBmT007H1vRL1Nnvs
WpwJjycqXKNdMCMt+Apb6wXKeAFXhQJj4vrvpD1+2sWerd4wSnkBFBS2Jk5jO1k2
QXrlwoJIs7mTetaogLYNYuzSkrbtKijg9Uvv21+r5E9Ei9wENzIFvwgsetMhGtLf
grFumXEwtLphfV7Xl4P1bmh2xQJtYlPPRMZ+BEyR3EDkznwx6VSZuNmIaR1BHTsb
uKpP/CAgHEYFC6ngFXjqqcI3rq+v1xdRAExeCJppLiSSO+hp4MKXak9RjSKzFLw9
HYEnDQAGzKy7WSzEO+gCs54BTTf6YhJWalDZFw39o0DMBjIHbcwMoAUQXq+IYewT
VvUoKq8rfo1uiNm7XCZZZJlqifkwYHWBZMNCC8a50TLZk+6abekP/2nkciVJIaZG
o7oIN5ZwPCaXLsie9A8W/DJR72r4wv5Zt7oIn4ZALgKtvNMn7iJwC5lJRkeokULa
T61/ranEROxulMeY/uH3FQcZUEELdG57RItXnnJWUFiFw3W9QAQ4Z7wRXIoheOYC
eMOCN/DO5ruNFegDDY3Mq1h4N8K8GUwej1dTfAUDoYpm2LRE4d5PvjJF81rOZlqt
TKy51J0nDrff0bNBAMdLu19AgxrJDsNYNc+jNB7W9XZK/WTJP+crldoy+7uuRx8x
I6gCNT6gQq7evbyjnEh5Xv4P7AB1B5uIZqmA3dJl+VXjCwq9Fq2huj7hI/1yp4qs
3nHKDsOv83P7XXrNsWIYSw==
`protect END_PROTECTED
