`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePD2/uakF03JVrl8nrKA0ApDBzhs7OL43wYKPTNL67nz
FxAD3eGdghHNhGX091uwfNRFlZJ2GgmgXbS07mxe3ES1jCl8Q9J/rmHd6cvFeBec
uGOqvwwuCfJqsFfWQeBV7ToWIfL23/OmiWapqxJNSuPMlVe6wUcibqe2pDHA/1Qo
NmhgRsgHvaNNa7853FcydCJKxpdHXdmilOU0SoFheln0mSn5DSkxJ3MFpWvnft20
D57cjP4X7x3bCiqx4ZhUKQDolNUIUIJexb84xCSyePcgt3RrRXI77OmwAQVjugy+
shZ9kZcH0wX/p5r1lX+IERvJU509Lp4J6l2foFafv+m1N1ZISICHnzMtFzQ/byD2
3Ia5HH3HZMAxNoPuuFzpUD2dt5kaKpAGpePyo5BwgCKPzy9YdygJ41lm4XkYiM3K
cTipadQ9UjMf7m1LCAXKQug/6+q6EX8gPwXDe0SRYoFeszlfaOny8oKjxFYbRPBF
2mkMevWoqC5PIn9TSzPgrPTNCll5ahC1eBDBdw/N1Ihuazrij711MFwlDnF6llf/
`protect END_PROTECTED
