`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMLgHgx0XXu+H0a5QidQl24z4AbI/s1RGE5ROzGlTu+w
dV1cbJeHHONSEovdlDeghzw4pgFK+Ev8dKRyauQGSBm6Nj2O2uxZnsppZ+TFh0Ri
IdQe98i/3iaA6t/pbPk9xE58FZsAdHjSn+TMRvCh6dj+T/AT2PE9Jt7gFiiXBavy
0TIApzXjPT9FYBPeDJVEPg==
`protect END_PROTECTED
