`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+Hon4PDnBig/3mYOiBL62S7uxDrvLJNsgm79jz95/Ef+ctlZtw/q51DaHiR0SkIH
OR1WsXHJinn5Vznqm8s4mWgphLtsznokzHDMBgd85NuR/lBv5wdYUwYWhguHk4Gn
rWOxJ/SAI10fuSzwHMcvkhuQu5xP1WbDCtQRh2laV8LXoBY+KLK8cuOq+KgKze2L
bkmg3fbCKwN2/4xF8KZTxQXv3tZGL6YNGjC7hu4tF4U=
`protect END_PROTECTED
