`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFYo9vfR60Gd3yE9m/m8nqV8zGrxg6WtsRjA+wWCdlwS
EcbUtYMeEnsdPrvU5gyorO014tV2SmMUUzURg3vGoBTuElttU+puCdRcwc9LmopO
8/FXbMG+dqkDP+DKQ5f4O9YFqmeiF9mfDfeLjAUzjZOHcpfmwYHuz/oeiM4PoITH
C/EYkB9Tr8MNzbNBzopCOMI4cI3B2EExplZOrcfUtOU=
`protect END_PROTECTED
