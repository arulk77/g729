`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL84yO0mxGno0SmFTAnQFKgcZpVdGNDaEG/SfU6erRmcH4
u3OXRNAZ7KTw5Ftwc2BZX3JMHDSe4MVliUza0ApmXxMsKzCGDeo1VroSGXlby4EM
rVvus/gJj1e3fVMfP/REtl0y8C+ALkRtzm3CVoWNro3TSHbyOHIhZm+yeVoRLZJ6
T3C5ZUOoyVnhl6DISoAhZ4RYneb/uG3UyjVPMWUx8EUg3uZjZB1Clz5Fs79i83IF
WWwYQnb8bTBKzwX+BYZ1h5q1sCv5JpJfuvNRaKKjizRy1NboPrkxd96rrB/1j4Ps
vnI049qyyA+WucsbFr5+QWKfRjMcBCruJNi3+1X+BzFEuKbwSOwWph5VaT0FKjwU
RhpaYhiIODpY1PUBaasQyRbf7clAO7cX7rRdX8k8XIg4jer32uxW0S3I+ztlwhzv
zxM5JCnplCf4Dhs1+zCY3Sf/tb1mUTqKyGNoWTqSQXfZTL2fyFU9t31EE3YdR1iH
aRjZbyDVJDwCQ2zt1Abh8kJvzwKOe+8FIbPy2oVapt4nfWGrf2bV+dp4SSnVXVUw
cFmE/deW0zmesi5GcVtQGVwCmgVp5Nh6Wecjo9ZeDeGvVd6chVjQ8IOghu/p1Gho
fDztQTG/2lW5mKbpg/aUwnQYEmFiowPBC3AgBeckGPzRGqexL5AzWZ5Q2NRUelxx
8Mg0Z83Psgv2ztoX6JGuA+zkqQynVr3NP8VO4e8RXddp2RPSWy+WGeQlXGSIIlHH
RPppVYAgPYPL+aTQnGUPpW8XxBLKsnDUC6JHUYZYLpQvXkwHt/SL4MRx6X5bJ1WG
IS+r0brAeTxgn2AMYLcwe/RazX1kBp4HMfGbJJRWtfw/RnX2NgPuAce65bAEX1vA
pTuE4J+DdJlZTfajfGn91vSuOKo+5ZVChzDqAhXTG8nFo2YABpoJD/2ww6PB90P8
VP/WZ/lzk3nHarqv/nvrt5cQ0jJ7iASUxb94MRYQ6PrUy+yUUvDFOY0pwj4Erwqc
WP0NDb/0ZzbJO6RS/qCvi2ny+685QF28CHeYPfsbJ7T9mHWWP6d1L9OiJWV+5x+X
`protect END_PROTECTED
