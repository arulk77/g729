`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4y1sh9JatrPUXH/ek/F5l42nuLIE7O/Z4fWQK9Qum7qM
yeNXxJ4zx4NNpSvWg8/QCYh8/Y8zkOj6OhWKGSyKi9eWtkW0c/Gg0oEg6/ZbO6/J
e+mtPjv8JeiZHO3bYlqIKEEMzIoSRMdPSYoj0enY3glyRJO+wPKYRzCwueS8M8Z1
a3LAuNqwnHqdRGLx97eVJ039GsfQw5dX5Gntn1WehP6vPYDOc/KbI/AweOTMcMjF
qY2kW7bgk34BnGrm5aAmqO90sthDDN3QGiaSO8vcED39nV3+FmNiLb7XjLGQtzS5
g+vKBCIB+oQSKcpJ+dZ5IvRAwd/dF+tujTTieYSJEfk+1/xzt0DZzBfuWvryLVjp
YfrHei1J4uzOeu7DgBrhaA==
`protect END_PROTECTED
