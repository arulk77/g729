`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKBa9oM4Kz/8/NoJ70Dp//b31eSdIFYTn13PuAi0JWHe
TjiY75lD1uMZYhkX9CVvpQK2GkpYPYUcW9v4oqt1G6GPc2+zgerpo2HBtAysuiq6
tmcqAjRb0MXOi2XPzoDZIJ978WTud9r5pFXdo3qigsXvT2quGW8j43m9b4mshTdV
/adGCQ2bdfcWE+U8Q06i6LdV+EwSd9NjoOYUlvyGoS5E0Yyz32+95S6of7E5AzRN
P2o2jUWQsReON3cm+RjxY4xNvNCUlmlQ1RCZciMjW9sOc+bLVx3ar32+f3RuyOT0
K3YTQ9YQN5zqKhqRbe8LQ4u6gifnVNmaUGL+htRUUqnAxjlmO49Qf6jZEABYumlo
bfuAGxk5t6DCztMmyz96wDrxq2ER0zBVvWpP4cA64sX3K4v7pcSYa9GuBK9W2+li
gkHeYkRm3CF4BjN8lp8OTbW9OIb/TlzwBiUpFEPB9eUbgm1qL86Ga0GtsTRRDFuZ
ZSBgONMELh3e3AfoQbN3/Ydn9SnLDY7pO7j+MSIAAGGJjVdx/oql4Vq7CUKeHvoO
`protect END_PROTECTED
