`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu441K+QVNWyjlsVXeR2oD94tZP+vQpxZpNdEU+xgszLB6
SkQqH5UtU3uipZF/6VVKPT0BFd+/a+xvp2lQJDOzK4sog5BYhEp5wADzsM98wTru
Gj4EW/5OebtQOKSYBBXGEidimKgXN6MPq4P1+wz2wfL7P5IpyhjJp9BpSTc3C5wr
jhNBqhLejP8noDVQo/ua7MzME+xR7biUcDq80gFmmHVC4Cico3XZgCu4l0zp5S8R
HehJlhiQ5W8qfZCBANjR07RaUO/WsUxp84MKNDEr2xxAMP3wJyaTQGFxoF1UeRcP
c9NuMXYngcLz5hca6HqN2g==
`protect END_PROTECTED
