`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJjLrOu9gQbStpqmmVF3cabRdQeeljS5rmWLpItL0d8c
gyeoLPQc0CHNZ6E63Z0mNo+F8YqEH0PTi+G9cYgplLSMDJzwOFB9QqA2hp2Tcife
bSN580r7x+9nw7oMSRK0bLzY1skl42TAQLVwoVHOUBz1ZV4tQhww6Q0Ookvs66bP
tNFP0vgPo3XTqbDMEduNcb/IdeSg+Wcho3E1M1ZHCKe9tvrDNfSeSrsqEEINEU1t
`protect END_PROTECTED
