`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGNl8tXZCHgVy9mKdy4KMT40sQP/wNb8qgigLf/LNSji
4xBEOJx+UVgXd974N/9xZoYRzNj3qeDgwhPDvRKJz9p5iCSW6d/z5GaS7MpcI2v0
bONmeWrKiqXiIPjKs8TTNPz+LB2COmpHQblkCxjVY3MPXX3Rcct1qrVvKMuoQyc9
ztZpVpbtSegSEJCdu3jtTaAJ4UmB0MlXXDyuptTYClxcIHJP86Hdzez6zNuGvcPf
VrkhHEu7ReSwqG6C6Nj9/VibMEFOTO7Q66llQjAFF+oT/uWgVvCJZxfYdGtsW/OY
GXTPoUaX3ILcX0WcUuDGd6XulkeNL//NBnxP/jOrITL0AY8Kit3oakTmjgfgrYT2
pBfXp++u55mPGsrjpzcrSi7pk5hqjAlLj5+R4faZLNmr56SXpn97zMKOEIn7j4fI
PVP8QYbqDMIHPdwm8NQkUC1t0in/La8Z79rZMnADc6jj3pHJ7ytUFM6etcveX544
EtIOh71mcr8h0rvuG6NL+IqfmGqbcqm7Z3Q6qB4RPMk=
`protect END_PROTECTED
