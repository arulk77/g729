`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFxSsx33qnRoZIJxdjaZ6dezDZpQ93x75fWtxZxt6EoL
vD4nNvFeFfqnIJK6rUUdTgnc97WVnWK8+YWpejKr4eMA93sSvPqT4MxiheBjak+p
wv/YuRYnomCY6la9kpMjKor+btC1GjbT0tL1jmJWKWPpZsHC4Az8bBD3l6Xw3SB1
bDpl/MChHG4eBkY5s6ZY/FF2+HHmhr6unf01QyP7Qy6JK6zpQ7n/MqqvKScPeQaX
mBALRbn8mRiBfUL8ys+egAX2ndzS8GvbnhNt8YvuxVFh7RZHkVPqLpebSjmcqBES
OcGbmkETWp8T4EXhGRURHQzqJ2yIGy4WL6i3GAZehH6YkueFZMoNBqnNRX8zn5lT
MbaWO9psWENJCC2d5cGYYJG3bv6uJzfEEKN1ONWoJLb5OjRr0ZhwgEf+OsxPMuZD
yWBVVC4CHlK3koKCjN1kC221+zv4fROWlGv70Ws4IXNOmaDxeHO8N8+Xpm+LvBMR
uxoGKbwVOj/0w/bf/i2URUtFH9GlOklQISQNsbp1s9G8jwWCEBgNoGVWVcYCurN7
`protect END_PROTECTED
