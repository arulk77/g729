`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Y2crHvBg9YfrbVEvJX1kPnw2Gfr+atj5uviCT/VDHeAYOvNp3ZC1jiIM3bY33uun
CD9IDBrpaUMzZocv20jFoRW9AUORY+i8ua5QL+wN7wem+5mFboQNIa5tj3rVfpRZ
2FFGHj4ONrrW5128TDYeB6BStAhKGb6koOiX3BXbFUYd+H+fqWMJZ1XERmgsirCz
AlG9PiMF5sSKzrgrWXZBIHuyGVbRlki1Zse2a3h00D7JtjIvTwaYsGhPMLPqYT5N
6/VVBU8A/miBA4HZq0mSOrjMbFsbV91gSoFhW5PotO4=
`protect END_PROTECTED
