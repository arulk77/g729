`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
w51KVXYAXknMLtPLjrjQEgOBMuBTSzGzse89P/1Bg4qso4KWrKwoFGUHDUAJaJzk
dBecguN/uLeVkrCT/4stIOOL1fB1AzqJdR64PIBWyIiRQuolmc4wYFaB4Mzt/jZZ
`protect END_PROTECTED
