`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
heo9ZRDzWNOi1gFAxWiva1lE7XC9t8dIonBj1orrW+JYD1zKr2DFPOHc6QPU4qld
HhQV3rgKkiP9UM83HTBgJrsgpdv79Ny7rw7nmbnXXU2ijK1s+3gxhnsll/V5C9v3
/99XlUc0pY1IqJMCxdtzTEuwl/t7ReRa+CsM/VKwk5tvBQkR5Gtvac+N/YxCaMjF
yX6CfBd9DtQouWJuPpeWVAT+/ETvxhUT7HqEzuvh/5/fcwfHzk+j4s5F1AeF0x18
cSzLICqMvwA0SMV8w2NZ9bBVRipxLCBgRCvk1NwJ8pNWCHwwRL8yjpn3KqW4BwqI
s8Lwxuc337F6cpuqTTCKI2bPaRP6iOo+bf0Juzb8oN2v0/rDbISIdBFj2R3omVlE
9Puy4bwEWDN+Rw5N34l3sdJAFOu8gJ6F1iIzTgSC6yNz0Dxs7/33bAcKqLcX+Jp+
q1OEnpGnu5SarbChyg7upFYaaWmziP+cpHNqAHlzhiUw5Qj8gvgED8/3oYN8DCtr
jpG3TOu1Au7pwcUVmNPfQSuAbT2j8KdAAy0FMqpzTghHQ6Xy9whv+S3H08nYSneB
itB/b74ELL/j6kRSdNRD4bHQ/4Z4gKi4cKsC3AK8AKjYKGpjXOcseHLC83z/EE1K
2DvulRc8bokNsJP71WQkgObyUIKVDIWTMDxQqjAJw5JnZaseY19HrLU7yrslTleP
HHmq8jMOT/ZnDEIA+/KZjXeF2BITkSL4u0NIAhNKrNuX7/mYMlzCxeiWaReZReHp
2yxLBTK3nRmrR+Lq7pNTkTa6pqTNaSEDAtd3g4lwfL4p5vv21k2r3Ocuod+O0BNS
j73AwjO2sQ/fzlEKO6wWa4AQ5J1rwDNNpzvL6mpq/GxP7DLTFd+wsxLMUmoCTRsa
UmSvEz3bzZflp8LcmaeMbqxBsWWg3pkjte79eIyEsIGcatxbMZ780HUpTfR9ke5v
RHSkfRJgtxgB5TN34v6Qa3QeMpDs7kDiT8PvicF4fRZaRdk67GqM1J6OWYbB5MGP
cUbYtcXl/UBU9sXWsxcDPWBYrVd8/DefqujjrxGnPhLQcUcbNCFAEqhaZyyxVi6K
zNGMpHudN9/YtLa3eP6wMdgeESKS2j6v6ULrhRC+hl/luijMTOeHgb4kfXt7ZHss
ZORoblxxuPnOLHyNx8omtQ==
`protect END_PROTECTED
