`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44fVSER9zXZoMxgky50ziMjBINq6xW1G4WNQH0CqkT8+
68Q6yJSMHWrzOACmsoXTYMHAJ43Wwg80Cm7llIEnGbibBOrnbj0wtuK7Z9UPCR6Q
aOEASCAu+nJ5ynkO6QHHMKnEoVMYfJMzWFXX+YZ7O2YOCYmxFE2wi0V40kGQe3rs
VtKSHAFxpvyfN8UHz3V6HPMH0Zeh0PFojZIDWtrSL/Yyj7zC4YLCLQljXXtWUaM+
/FimCCCSM19JxC//hByNpVNHGBynZTo1wP42WXJ1fuysqnUUyta9hnZP22K87z3X
ZBbfYhMeIAI25IsCKHezKwtsDetLr2e5A2d8W3Yfp9+shUAIHfXRoIjW4IuIuQjD
ma/BC1bl27KYJg7Nz+gc8w==
`protect END_PROTECTED
