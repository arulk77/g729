`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abusY2hyZx52aAUFeJveFHQ3qxc419jqZReAr4PtJ+mO
Ic0YiXijvSgu+i33aC4ytjthgg0fJjtMgv3eh9Fhdz8aKcMcOed3mvfaLmlilIg4
kzn94UyDrXHZkZSXwYJlc4ibn87dgdt3run8xMji8l7OXAficvvlPbp3XZj1BbwP
Txq6SezXXEoriTkPuAiXJCJnBJMqhGn0oGpURiEHRdrt1ef+dnGzJQOu33fWDj6D
xrw6pDN8keNX8/waDoML4yjiGV1fbnDmLeqX3gnBi+KGgDPp+xvqVvwk1fk1Sn3X
OBekBnPAUIMBRJuz+vRnB4dSGVaAuyDZ97o/CjjsyTjwRv7R8BQgK/82y+5qqR7z
PN7zXZtAQERNe1eL90jcZwJDWEvuZnWsXY40w34b7xHRI3UTF34wi4qDZXdW8TD7
SsYgCP0PE41P7N1vaKAopwACyRiCk3QHTalVEhXaJLTJQdnbgYjo0r15jXMFMnF7
cBi5GyEJb01FqA726kOeY0i4aUPGPNJcQzyCJEyUpUUTC2MleV8ZEuOVwKExD+59
2e+R+/zTPeZBwBv0iVGbsHf2+0AMeWl813D9VbbeoM4MnEqUfbqaNOaIEuMrbkW9
TrjhDHIAFxa20VY9cBDJCSEhmEUSA/8Gs0nQkZJdosyxdQxEj9fhaStf4NA59kwS
/sV+9RAAMXPvoBpM3lzy8JvBJdi/Gb4Gf+KoczdcL7xCCRjez9AKK50+3h/n6rdP
Fd7KH6xUnmsOhrLsWFUCXlDWriM4vqy19abSwkl2pNU7dNE6okGuzVoGn0/gDRhS
dJTkMwarYSZfbFUKTuPjnxf8tUFMtqz62vBhhL1vTIiEZJdUyoEdkeeqKSRusm1U
c8ANyIov6BkI6kqchPMOzaGGgFRCm9BBqmJKZYwhbkgO0xoJ6kIWRCQDVXTntydV
PU5BGxJT5DFFsU2C/v/3RUK19myHSxp+FaAxCaASPqpUhKdgp5/5PBggzlXJwPW6
KPm+xHucaBTv3oD0d41J03yN9vZmCI0PJdXXGicJ6s5iW5G455j9QO4iFfu8rsf5
EU6wTu9ZxfR90VAouW2bmieIpUaS00v+Okpja8zT6EqhH7pPyWOac/HXNIzuUFYm
giT+TqhpTiaCN9KSAASk/ugegLZgUePG3OdvG4zz3p0dV6FFkHVEpB7ha+UPaODM
XStZ98BV1bXfEkB9FDTR7Uh986wFLzwQXPDgcbqlruE1XEgXvVtsNioOim0K4Z9R
anT/bk8sQT/meFUXhKXPOAOzVkQhkDPn6/fu/TDJbgWI2pZVf7gLmvKEP/cw7vFX
DUU/rn0qZBbqArvPQDfTYqaeVldbq5pjw/kCf6KR1SC36OHvccPcDvM8dLRYWejB
Xs6sqegx/8WRowAmrx+wHhu41gw6IZjxkyOdj6QXwDohpvZak6HUhNsF6juEDn7i
BsqI10YFGM9DmzvESoJqp2r4Z0NQv2vBRKS7xn9U0UfAWwUCw8V20g7VkTyvnj3A
S1TD0MaqGZxGkpfpaGbZQ+Tg7iuS4NKRbd3VqQPSB0HJARq25HmsQdFcMVll2cYs
l+WCPrIuTB63v/DT8FfSzaicXvCeWm406YWHHNoerWljx039RuxxAzLB1owlBgZw
COP8wkaRAI/OaU3C0EqxR/5+enKcYlyvK3jdQj4nZ59h3ey4tWRhs0zGJKP+HVta
HrrF9jIf2RkTURChIuTxqDoB64lqOjQgxbb1hkRHk9wrSyPHuDrNWVXKGEydDv9p
9B+V3PrXT5lMxTSZQ5taU2T6QCaiMTVagc1Kq5ey09lZhN+P6OrZw1OpliSjvjG9
L1U+bexUMq9gPWTEvkgr0osWB3Uzpj4PscM2KYiVRx4o7DtAnwlhU7T+xuiyfrMO
9Nxz3aVZfFYfxFNZPBSOGte9JcsBVeBR4J8SzzAIkVBhigASmLH7iggZuXH03mgn
633c8Dz8dQyel4ORaNnXi+IB7zyGgQcNH5psRzmkaVndZxJnQQM0/+FPOraLrQkP
7nzvxksQrlSeQ92fRoJhVjUull7oHnu57tviX9N5TXm1qsSmjTKa/1N6AfOmvbgm
C2KFQ1qEumsdCgyRtgi3Ocy3Ve3KxZ+mvWah/fSyQXD07e8I9yYgbQGSIeOch6K2
Ue5xCH19RskLs7yUFLaOxZaF+iDPtcXR8dMHhOD6gPWLVCr4onOfZQgAus5Hymvl
A8l7y8whRjwvrAiQP/C9CC5ofdWSu/m10IEEaWXTUIA6cJZF9hOQo4O0Ws/07tcV
FxakguTnRhugGpA+js/Hsg+SvyBqM7mlGq52MlPIrnLcKAvKGJRY0SGb26brQQdW
slAP1VGA/INrbzW7eVLCcsU/JdfBa+t/XIqAa9fMOshJGFsHcSXmDSnFwt2KEnVi
LhGGZ5st28NFtd3GZ8pd+yW+kqaUIEOkAZ7KQaM1i0t6SIw+7n1pn6Z8kzi2PJkc
DV0MsSSqR4xrCc3dMDG7f2YKvNPjb1nBc6B3ZD/2RRXMmFg4bv+34BjGSSSbIEnc
bJL2qbYSxY+nAvIEOb35hHWRRxJHYtMWPb42/Oje3o+z6WgoSG0NM1MxKCqAJlTX
ulJlHkCuglvCYDWFHfLfD96dYhx6uDkehsmPXJB6KXdOWmyPw2vRSsabKhmonm1i
F8X4GO4VzCDFrUtijBARmsfFqb3yVgfGQpCA1gmbjTh0iIp/PPZPY7CIGsfpbpX6
OJDtkO1h/h/nSQAX94uw6kjnKgOy7FyyGzYxTsfSFgqDctRFt/chbbSwHd1sFWxe
Ah83iHozGmRpJjoeNpfIaUtk5n8AbSzZRIfUKjCzT5pM/B6TAs0nvtR8e+92LtUC
D9waTHugb7IR+ixHt2Jc/TVp8DggTgV0d/YWMZAhx6TKO2tMpvkNe9YWsKbCiwI6
Is63HRSb91fFfgQVfX88y97lA6wpf84PQTMS/5j0yI1tdva1iGNRVAwh/XzePlbq
QmaqQhI38KKozhnoS3xVFEn6CpdvkC5aXrr43NETPlusuRprNvG8ejonrlcpTdx7
rbHh4qbUa+yFhUQRGLaqh+i3gCrlKL4Xa9u6EJrHUtcMq3PwlQT+7C+RZwWZmEVK
RLcz0QihFeVGkk6hX/tntvqSej7ZX4BxSsdJA1xmTumF54JdWNCyj7NUObPGuMJc
fousx5xamh2vL/1gXRhSMg223mDsQV6gbP17Xiqq0J03LINhtZkqOOLl/1l+O7pU
+P8cjuotkQUA6kdnD8Eb+Bx5rok/YrN09e9WMvup0Ij5JQlP2vLKJ/03WfsXydBS
DQuPmCo5TqPcNzBtdZOqXfjjKLcVcN7I9UdD7zgTPLz5pnTbRRjHfAmtltq8ujJJ
IBAMia7kCtIHwtQ7+XYnT9b7cICJEnK6PxlVoRS3BxTbQ7Af4ttGhzPquSn1RdmI
HU+7Z4qnhmGIvvJp4PLh42MkfdGIjqi+V8hx8Li6bAb27CaC1ns34y221uXh/twg
OFWIljqc6Uhm4cj8Rvk47vaQPli3llqKtKNZOEXVSHGDwV6w4NO4aI3HAsNMuoqZ
FaCqSl6vdtCAAHzb6WsQXzj6euEud1kQVjNsHuzSkBp4EBQs+XBDk7eKySZ3iDPL
ToIuQbhNRW4xsSRazJBzJyWUDUl5iOUPb9eN1YeZHYrMLf0h7BeEmRDD5zIbmA7j
4qryCXuor5NhzzRD40HXxRRm8GzWMjoIMyQtToAKqDwynGhlN4unZ3rC7y1KmXmR
/ahnmRKhrt7xy8nJZefuxEYa42h6p6WcW2xg+54oLjwiRL2uxEY5MvULgITNH/EO
Hptg+Rkob2whWvzxJGpF/C7blZnS53xfeZ1kXa6G2JF9w1ip/Bv5lKl8n3AqeP0W
OoCVUlpKa4WP3QpmgRn1kbDDisXM5pu+djBIvukhzn84cBrNs8l+HI3uBdjXuBae
LnQ5l9b03YwMRegSLblSMhnRnk5CmftK3QDBiZjwQEejeghbpYZD0fR+LSC24wdZ
sW7Ze32yxxoGU5+OF1Ix8u9NANndjMZqmPTLUIzq3Dilb6LFNZ5sGxnvFoeWFlmo
zNYjRNvWS9A15+WTdV72pJW7r1jMTx1eEFIAbVWLK/M/ttNXEsAAv7iBG3BpxaV7
K1wAYARiKLO1j4XHGUOXXuGS2gk46FITV8pAqYYg+m+DWhh5xOb0bS1T//u7B/QH
6cCG9rWo9+GkZVPnvCp9V1O2XYw8DQjn+eR6OkF9Bn0qxg4iSmdSG/47qhMAwgHs
LSXUoSu1b1sPo7MAIhxq4B6BOb8UqkLorkVoIziKjYWqZg+Ge7LpGkLZKYFRcEXs
mCN8e7dnT+vDibbzlxUE0V8vl5EZb2zcCcZnFJUq4w2aGVa+srg8e/VeNm7uRqOa
zUEel4cb165qx1n4YKZmzwcjjDFcDmmyMH8MIW/ef7d2tLUEGtpr5NvQJQfmbxFg
v060axjEo+9uL80Y1j8JjZY60zE1UYK1F9lTdvEQ1xcBCas7ROqFpjB8qhLcTZ8v
00wnsq9QHv3x6SjnfODL2UyyOzNQlG8cQ4LBNNnnJ/XXZwF3Hog7sjLAz3YzAXQg
LeWdlDpV/ajvLuJOnxZb76QlyJwx8w/NoClJpkmztVn4GgKZqUuSYZK4BbBOHMYP
oZxXI3YpHupKhVQLmOqFqmH47gNoetBL0yGAjuGGZE5m8sVbUn0b3ZaOgpM/HCgg
CWjCw8PmFmCwH3W4G6Nluuew173fYze2+iLjjIkt8nQ5VPvhRucRoUS06oWv84Rk
rorxs6Ev3yucgROOpu+Lw1qDzoVNknGBwhKd22gze/pXEF+TNm3LHPznlkp9eNFQ
8H4uhFN1/6B9203RwsdJsLUZXhQo1LstzFU9C9KPoOFFBeIk1H87YXtvNMmo36XW
IzUpw4q5VIF1syk5D+JdhvVRtCseirnlBXLDf8Pa/g8OvIqmDuSWhEGRN1TqZV9y
yjBSiacM9ATCIiCwJvKTGWujT+Mj0cXuAc8vUAUyxwjRminq9Ht/LrV+Fq4tFEp8
TXW5WElnyjaSYHiHfuXc05aiB8lafy80MXMFYh/GhvZGGYiFAvyxL8kYEBhMwF4A
1xScFSoLlYVADY44uus3nUChl58XWTb9NCQVKPzJ9FNfxe3DpEkzc3AqA/UGFBhH
JHn+Z+OlQqb7J8+ScVPiOLDbByMVhGnyoG3JsYNDV5inhLthzjm5g4MReu6Zndd4
LEjFZ5gm/v2wIxTgwdr/H8eo7jDakkK8qqhMhf1nQ3eeP0tUavFpKy98eAwV28+x
c9CVhi8WcAgU9p8RVHOHgjjYsHAaaRZZBNtRYBLYv4VJ7mlWUaIBbry6qIb/iEfa
OLoro6gKf860wKWvwAZbDfHlSqeTe+W51G6Msrf06T0=
`protect END_PROTECTED
