`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGaA85/mTuQj7m9BOoikWC1gVoHJgHNXh41jANstEKHI
nkx7MhU8+8fK0iBgtJVQ0/CHXLsPvjmRrcHWO+YSbmIWuX3I5TLt/RSYtUdnNkHT
QjeM2CkXJroBTbvYC/+oQMzLxurQFyGFfslNVtOTEEikINjDuFq4hyyzeh0DtAOZ
PEvc2HaOGdaqojClFU5PfM1pKz+fjcUlSX4BTe0Rf9FjLP+fmEnqVzRrpvL4ysZk
`protect END_PROTECTED
