`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SRvkL6jgWgEFEk/0wtk/gbUJL0nlZkBbmcIsYQ5YgDbI
FnvXEooFhaeMe/6cdmUhMeieENA4kvOAwLxWove6u1+ctviAPBDppcXXJKmqp98n
q6hTEstov5xgLpceeaJUD5uhIBErSbqecBljLuS28Aa543l4ozOnoYB4POmg5bOZ
OkS/HYcN+K6sOQyahK+zlf5rK3nM0QywsZS/8ke6QDiW2klzbrKo5RW4OwvvLP7t
Y3MDeRlKdIrvBK/2TQa1az+gHG6uPx3LLrmAlMkc0m1MeazNrZKwoUWJOBnpKxyQ
grWY0+F3m9GbYvOgjyUyQ+Eeq0RzqcnKfA4Ki3xrtxZLTkpbhGiCSLeK+A5T11zT
38WccGluCfZ7je3C2UE0mHyV7wiw2qYllZLLrZ+SnC5fnRjUDysGGCVpYMhbbhDK
+UfnIh3Ikhm8fgaMtwTtU3Om+pKJe+lqtX2hmoAbLL9Wd3Q/+RfcCNYq2qH5xDqH
xci3PUVfbwUsPro7qjAnpdqRVqbXMqU5CaD8qkIZO8t6YOR8MdtH/exC5lSiAu+D
g9RucQ3lz1Q2F7K1QXuoNzfakzRXxZF6Y+nlT//Z+LY2rXs/HBFoCFZRzw3SXiux
AXBM7HArm7leOr14WBHfYKnrUTYVccGCtnUFyAxxUaXt+caiHtTfOgU6UbMOolKW
lFRKoAUGzYMtHq/1QHGmw5HOtIK+dLZOeVXRXOGHeA/4giS2h7yWtgBMe7xde8UX
B1iyQqr0vPEWqmBh0aehKILYpiduYkEgAQ/TCbvbWE/WoMvuv4RAIPQv8uSattZ5
G5AWJgQMF7MJnndtj36iWHeEcp47O4XCMoGFtcIW2wOFeP/gRrZb3dh6zrk9nfBi
wWMZ4h4QCfknQK+ddw/oxm1tRynVJTxctBGSkZjY22zE3dd1B9gq/TxNXaZKYuVe
Tvov3i5oJRufK2kfo/OCcPU2d+iKLCaTnp2Ktv78CBx+ZGdBIcPhwmIFI/mTOILl
Ce6YKp7P5dpPT+7PJykq/e4nr8gO3BBiO7e4X9KwM6YSJXFzeGM99VU0l67MfSaG
2zjxZNqjiMesem8uMeKVMsvEE4nebswRd0dqi96b8S+VreP481KDLHvmncFIoYVv
BhSzPYddo1XFalvLT7NQRMDyqV+ZeqGBw96okHuJtIv43U2uPEETtLjhyZQB3kvJ
t7K+07jOGwFu+vdZoGBD0UaendHoCsSy4KptK0QZ26fY3U4acqGMOB++Kzrc4ws/
qS36o2U8/Lx2fdj2eExJY9hC2OgXgcwCmfW4uHbeJJhKwAaOcsvHx0lfhO9fe7DB
Mhs2uMdyyNc/EfJPtNTS9mkGX6kzxz6lyk64/sRMol7CivSunMkPbAIt3ZpUdc/q
PnKQ4aWvbHVmd4x75s/wRBOqk3HucoZikvbZIzdLWJKq5hZ8uiFT2e6mGTM2rpL4
9jTnbGbvtl42/6ZWLg27ufU56ciCYyb1f2/xJ+EjtiWfEWmrTQPzmfGCqqITSmNd
HePFY1MjYfesr+PkaelBBKK48/VQ79c1p1fsyXBMkWqXmI+aTWpVGfSCz4cNoIBH
y7hobTb2N9o6czt145y7rbilffy8/Qf7xB3YDuWfhtRCqW4oCR1hCL4Q545TDAlG
eW18uOM1XRBkYhbalOGFPQxIEqyaz034hRr86AraNeO1voVzfVFtuHNyrpW05upR
IgSiQ8jdeci0UfHlsBpap00lNHABtdWI37mleyAdxNA=
`protect END_PROTECTED
