`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eQjoFJDQlr6OmoMjzKIA3Q0N8IufLjUZwtsXTLaB8JB9xU0Bx5oMG378qM7DoTeh
n0Ar+Pd1NscUqtLlwDdqH7cpWG98Uw85JGhYnTMvKpZ6gfnL8NJr7XVnYCfqhk4P
8vjwwUSstTZ/oqB9oGm0dAwK2prfGBMKWTi7Q8E2BiQvPKi23i8arM9sK/R9nxV2
ReD5I9My7er3x9SJ6U5vjpPhcu5za3h1wKdCE0NYa8IPAahLs8eVeamGns7fhUKu
1Pvhf+8aiWZbh7Zihw24urmgu5FWB7CdWpO5MNGdSIVpENql3G5yoAzvMryeOy+s
OttNCKS9WgG6lrJoVZ87Tg1ldap/DS6TF9be03BWpM+9vfYqDcuHXwsN4tgcVlBU
exEUdr8dmWj2zcYk5dxfuOo6iQVLTca1vKQgPF1Jn/Jztzbxr4zeZEdhBB05WJvA
g0PQ7TmfIAwWOJQXvQizB1LyGQR0mjGd6A5/6yJbIdTmDp9VQEQHrvDpb3XfpO59
fPex7rUl258675VvVMOgUQ==
`protect END_PROTECTED
