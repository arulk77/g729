`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxLxMs1WxDr/V5P+zQLvAChQ3r1JKxsjcvchLZJ9OqUs
KzmLwmhWy3Gs+Kg+QDHaVmnW62hgFekfECCAUZmuZla9DhVBZm1foYAYSgERsLj7
OoWzOTYrWET7GLZjzMhwpZ4OZKX36qK3N2fqCdWybFwgH5bWggFGwUy7F75vZyBr
o37Sg1GtUoc8ruSO2YD083pdLhmPrD+gJiJPOzw4TzFDfehyW9jWy9tRcOtS9UU8
h0p9GG8MtY2pQwR8nVa7XgjprrDG4Uu6o9Zw3xz7edGd7YkOOCLYoZG9FjUy+Cz2
BeABbTA5Z6qNFkKn3YY5p9bcDJKH0noK/+9CL0WZUgIBVHyKmBOopTnf597r5dsL
UWQn8BgbpFoIHdURuMKsvxVikhuWCFFI7ErSYwN+HcxsrsBbD6C8B4yAzbPFX2Wy
2DWhpK7+FU56ALp7pGL8vHfQADTBMc9nUrLMknj3j1gGmNV1BhdzdtM273O90p0W
Vg5w8di5kyRPmMMH/k+2R2yHjKw102pZ15Q5h+k+9JIg+mGFLKiKnxKYE7C41BVk
YYWrnIPFLi4hMrkjZzMMCGnwDnoWlGQ6u1KWxxZAlkfoPXGX/Pqa59q1Wrz3qs8d
W2XVvJaeY6iG/Us+y+QMYDB5FOLYJ2o7nenSPCV4DiTgPHsY4STv7JJY5oQMWHbQ
YOxcHdjTBPRHDbCuBWjdPd+2JmQeG9x/mFviLjbPi5CTu810SB6C2uLUEMhL74O7
1hcqjPQM6nC7XGZlXakOeEiIG+zz+YTwtaKzOcbfnjaocYknR20vUMFD8gOPEEq2
t0yzyzHH95OTfxybe0/73jUFTCh8OlGMqKdw3IfnTFtSbU2z7m3X+pUOsmuTCgbS
GKyYvtOx0OoSV8PV8gAFcuzoqhs6vp30/6HzJ4pAMt/9fB5mLJqDsZFELT/1w77w
uTF6zljFfvvIb9O9Guy45LNoS4UKlwQd8rRlnRq0ea0TPOyWPXuSZOdglMmd3pjM
K4RVGEwORrqjE0hc1H52kTo0a9YXVZJogaRULK0YePv3gziQ5Dt9ewT5+8iHPSSR
FyLSzrVYUsmY9UtQzlqfTOXrtfR9Q5f68dF+U0ZGQYKFy1eJJWcexNJ9cvbZmI2U
fFL4OWRNRzuGyEO5yAVDwljz5IEr2WdvWnBxOxUiFVI3VmvaQN/NmNDgVOu8dPCU
zuX3ejQ7Fl40u3x86PceNGj4gxHSLr/XuYi/1hNOqIs8RpHmdtTdKK6mCwxAS5+L
zL3joOtlALNpy00BpiADgiV6N7tMjV+221RwDn9WP7dSWuk6ClXFFPNXni8kZWT1
+wLjaz9RWm3wZ3AEDg6Nk9wOznBoEgwU5w/P5tthU/dr0t9zR3Poqu6DRw9khOKk
39R3MuwLdiYaUaXKDw0PD5N3m0mT+SP8/lQFqIjcHDKwK39TuZt09hdKo733iRMf
imPLHQQOuMEe2Q0qOlY8ZNZlKexvzPJPb4g6ffcxDmvdS2ORmxmNkTeGTXhCMxqZ
4kWS7tHzR3TqCSPmdRdII/JIxefuQQYiKSve+1JqtQt693dfJZIl8xCHeA5W157V
X6WixmNjBFceZiLneZDVuvfAdQgkqxrVuZ9+8ZCOG6wqnBbfczVyQIaV5dmDIRYe
haE3XvvVpU4VD1ruqNNj4sPMF6MW6JObWh2IxeKLVRts4/VgGlhbEPIDI16fufrH
wDD6hSNeQdbHhdVaMA5a724drk0suzventGdNQLQ+SdCLjWx/+o5DPkOa7T8Jz7P
JJj10YVO0NFPSBXkRrhcsKgxjKWm5u7u5QkZLqi+qWuMwV1LWImk61cpMWNXFYMc
CYGE9u/BXE88mUDVtvzNWG0TT6WgOys4dfjr77h2MWnORU8PMfW6dxm3BS4BQYHl
ezmcu5I2RbJRBH8eyOwoqaVcUnw4I3mPnljmaJ1s4hwUZi7XlFSrS0rn7a50qTlc
n0xK0uhUwPgOqkcTXpWszfMKZ+FHh/GRhypqRf22V66+nh4LRBOCvoWYZDpdkCwL
u6aIce77BTLsJH9ZufUhOfHS1mehW0QJ+3bx6UvW9eSSO+iun0uPENANze4jSR7I
clkyUOI5o/WzLianCFCR+kQz2AkH0jTpd0CKU3HcYRVDzuC7W/jwCdLkck74FLSW
MrXoethFedPw7Xab2zE/G8fooFP/erVlI6QBUAX5KJUir43A+nUoyLfnlgwaLOkA
b5GmE0Ao5SdQXMfQZg71ryxJqtJuSvG/Dlqso551vAcfXqYpLfBpEilZveQ9JdI5
GaArTeRAykOd8tTXDfvlPTOR4aStI8er3H1aCa0yaPCY135Co0UoXMmVjNKTqoR/
92MtsTVzUnbK+3Bjzz1XpuWSWYpvb01B1faHydR0ph0Ditfm0VWRqxZoP1U37zSs
WczU1e+cb2Id8jItNAfT1qq0VyYXg02UqlRap5nGcL2ayCtlVIko/KwtPHqMbo3a
lor6QpB4YXKqDUivrzTHHz70+AJI3IR7KvWPMUadj/Rn2pVhOhggQ8raAPXe6g+S
MgMFdJ/ePgS1JVy89V6qiVCult8Bd+GI4iR5bkU1celoQksNjH5e+c88Wv+YgjZH
yGgMatxIQofSmMuz32B/8g5y4kzsHtzsiOWuS44FXDAwIBJeCPCwG1O3IkTx9ypN
E1uXw3Wzd/JrkL0pXv6q3Y2/0O6PVnguSgEkSUkZjUkqP/Nucdta6P9pyirBkF+j
Il5VJIY6p+oWiegm1C5EHdkmbN6npU5KWJyQzRDQ+OCgxzWo56tfcvx9KwWOCD+n
EmHO2zhBjctvXB8OJoc5O6hIdON3ndY9psJeU8BQvunbwY3YXywoI9W7y53G2xd3
PFxtNJ3AbNtQ5a6ohkRmWk1owboHF23HoLc/UEdk7N/MWZ1HPnRiuQKI0M8sRMN+
HLNg89FfZCjXuprbWe1agbFBbva5bMNjSParNl4hjV3xxE/4ca7fdRGxkQ+yECIy
SOuzYwamxvXhkw34tasVYJK0nLlAL50XAl82tf1qtj7fQiGE/8BwPR/nYPP/HJJC
mQLdiftMbYpEXqic4l+Y2So5O2Rjkw5tPZnlAnNlBIyxRvTAVA9CX4JVPGmujJxJ
pUo4XSOiXxnm4kkQz5Jxu0hmeXiNJFj4E2jCWPDNj7eyoS2CPQkvEmeSqtXldb3E
kR3byE0xY9mJ3UUrb4xqnUbxt1DK+K3tYMwgmTSaE+D5W0g29etX3wgLjTrDBlJ+
LXMUHxyOXbYwcdZng48VqsWuH8nodYt44ctx3/VVi1m5aEDn2TbLYemEGWueyJZU
AdCMJUDEuX04PLcb0lJPR3if1/EXutc6g3nTBamZp3Z8sq6qrfE2EQTo3vT/C3Ao
qMiGZBrhBUOuPiboxfCRJ0uM6dyPIrGF7XOxbAB7b3eUUtocVbdBAZKjPk5gamGQ
aAzEMkl5aUlUMvhM6B2U8UvkEzcIbI4PngPwZ5x5srjonAyzBl+jQ0yKRfbdLYnk
zGy0Mg01vrkK50XJ8AAYQN/kx3dZyfQZ/QTMrwa9oaUK8TahGiXKMN+wZG0Nm7s1
3NOE/x5VfiDcTiR2jXQ4jXSFgu0EzW3stoD70aXT2bQ7jGQA2lzIquZPttFKEk7T
U1KOglNZa8eV3HMtCIARIrbUQz3fHnTPKbAgZiwPP5XhwKT12qlLgE9wTRILFhel
pbS+YJ/jd90M97J9h3DlKXPLB6lzyvGbSUCwUP7S+VO9tUtEoZtu6Yl6qS033OWm
9qkNNDUqvunTbUdEOpg3T7FcUWRzyrQcc1hA0erzub08Ic254Mrv6Y3meNJt8x+T
c47qw+N+P/WYfX20HeBPRpJFkSLPU3u+ZGIzitrV4RkVj4Z92iDuPUD/LUHyrbEZ
ALROtAXvXZ9xStRux9PHzUXOdvzoc+sxO2+aMxQw7CPQWVeoRxxG+bRhjop4Nya4
DsMJKAEpPK/onl2ACxMmcTOGOY1vo4EtaDQJkTv4YC6pKVOtKcY4YstNBZHBPUoS
XLG/JknZjlxeeU5djGcOLSeuJVKD8Z+KbM1CF8w/Ooa3ci/J/b6d4/StwP0zSD08
BixJ1K8+b50dP/aqy5q3t6gvpCLPuE7kh3bSm1E2OQIb/KR/byowmJVN6Zh8EHDB
oUSjepB+d6f3L8FF7NAh5FCXjqdDN3HtQ97cS35PW2QWtCKi4SzE8f0Dz4v4qgVK
WAfUxPjTsjtZZqLo47oA884BCROW08gJDEQ0IjnazZPOaRIYDLQmfVH7u12kvDw4
RFHvHECxx9GXXQtTQcvP4GpMwHVRKBJH42db+vU8ADrfVYjaRMLIsyZ/u/ZkkA4E
NCMyQcstjWhQo7uj7QyGrZbTdP0FRh6yUoycnwugmxSWXIPqTPMKp26S9qEWujLm
IXxbQp3/riOJjxXxrlaKBBFZBfwnL9T0vmz+NdTmPPl/7i5zsmDVOZyN2BYTaio9
eg1YMmHm6+GhBZzbquRQUsb/IirAI7KcGtdTK2WdWzfZJKXPTCsVUPMc8oVeeLDv
eweTzKo9zbeqx5+Y+ViBpsAlWH+bhfRv8vEwyU8dUXa//zt5doOS8Q8yHQutO1wl
e8Ycxo0QhAzFg5zhmBvJhawaT9hvpLYrNYci8f8Tdf98I4WK7OdS1g3TrPzh6sa2
uzD01FNl+McnP1L/f/JzTaed34MjqEC+npOeAM/lnc/gn7AGUudNSLui+aieZaDj
GypvfVpl5neH4nn8QjKwtNZTMP7l1geqbZO4CDXA6ZgQfW8jEnTOF/Z7bGchQuuN
t/f+lXGUPg1ngPJhjB37O3lUUT5MdC2/1G590Q1hAa7esRGNf53ZbY0OA5PkHoAo
gH/XgwzgcJlFX/vUjwL9Zpz5qg1qvtbSisCl1ZfHFaOPJKN3c2iMFQREUf8cZSh9
3Fc/of6Mo8LNbuvb90+ROjh2yKeYziv2c0EY2iqYDVhFnsftmqBNVWRNf4SJHkEY
V18ws10mcH+CKF/wJVM1AJRLGTzxVeW95SMzb12VT4ylxBpp4hMnchaqn19anc3H
FVXqXah1jD2V7UllWXn+hjANUvlbAuDX2Bw6s1Ot68ajichFwp0ue4Ju73xAzKBH
AGJ2XtHeooLi69Qs44s0gmGLEpcO7rqBLbDekCUWgrdfCSSAOY854/7NzSygk6FY
gsMDjZNwuanGC0Zsb87LnHny3Fb/wnHbUV0SBhgX+P9QC336oyD8TVqDb39Mw+kC
cZeDkoyglrQBbQweP3Lm1ghQ1ripWARXRyyR7IyYoA3bqG6/kKfRm7sIIouvtXco
1jAF2D+UbKW6xo6xchWw6q6M0rT9XzCsgfVYGvv7ICLDtj21/rfFxZezl4yY+7gj
3AX6wuAIDWlNQDJU6a5BLY0Ja2d/ZfkbyRP4ZozXuJFpO/BVZWwrs1NnKJ7HQEJ4
wNz58qwyLRks+wlwmqwha+UlJfyApu6SRgcBj5ZM+QaggcBjQo9qdKAfqaImCa57
zLB5J08sSYZt1vF6SHE+Zho9dXG75OLxtpayqLCsiAYlQCpo1cKWG2J3qvbcwwVa
VXv7IOcQ1Z2tdjwldQLprckOGdvGCiXZot/mryYBZ3qJVtlG3oSCyisiVjVBTF53
c2TEq03GTKkbbaQKE2FPB9TIelqV/0tsggEtb9G3W/vuqwnZn6BxFGzsUk2vLWdK
/AcLnFUt9DC1TjCsItpDeX3anyWMJicatD9ZMhP9E0KkEJVGZ0m0vRzD/4TPG0bL
LpVkFxnm3U/AmUssfR9nhuB6R6ZwxT9T5djBaII0TCSq00pSeE1It4GdcS2m4ccH
i1mJe3aIgKHfREzgODh2c/sN4F9+j8cPo2Jp3RM2x03ZnC57ZiJBGKiCHCbC2hWW
bpK8K1X0ppzR93puKDcVx8ovfN20cvFULrehzON+Q6nlIgD7k4YqSOwduvEKbEGt
2bfcCVBPcevSiXabNrDsTZ+725DfT3QwWzJuz6d1FR0WN3R8YyS5uGWZaAfVU7c9
igr9sK9ywYi+6TomVWqG6yLs+vQL57cJ0Gm0CYkcnPpA5LnFHF7IITwNR1T+Hi23
jCIkoPAlWMvC85+LvSSMyrp6l8Awyt0qoYnYK5jswjUXarMe8kE0sqVvczu2lDwm
MbTsiF9cgS+aMnVhDd7hTC8x9Mforw/ce1OqElfV7zhPYLfIfgqh97RNsTokJO2d
OGiFK7idcRR+QTC9kuGrnmvQJC7BNAGx89yczT/NT3J13lvT4ymvmyLJF3JsQ/I5
qSlAc47sG75j9JoCkETFQnu2NFp4q2J/6jZBFUc2vyfXAbmRXB4O68PeITKsB5nG
OQQmkt2JXHNjIEnbFt955Bcee8BvmAS0fdhufCEaqN4GRgxtRwGgI9I5eXUm6Io0
hVL8KIu8Z52AFFIgES1Ou2S8n63pcVPu5bsy+rxtnliflbloMLXWVzMkiSHE7hI7
NJiwazbohC1/WlRB6OBOFczChcRMOCH3dUsD+4vOAttUHwmleEyZ0DCYdenAf2ax
niC9EHVVqZ0/i9XGUQzzKuOpZQDZvoSsHeVf+1xnKl2FRM2Ku2dt42A9h1XMyMJb
GuNsuypNBWFSWfYw64ozQ22RMRh+eX72SNqrqzDBIXcA8HDfTIpXvCGsLmMvPpr6
KFbzaD3ynEGLSPtYz8keJ/8l/IWYodysJNJtTlsE249G0ykixQJa62ZAeML7CxD7
gBTNiM4DqbWbLMdgdso3g/bsiiWakFmZSr+kxALZbqigYulPsh1XNywrHEjCZGzp
AovQXkoXIFjBM3hL+bRmYgh6GHfByyk1xvcBOi2MsdMYV10mqcDWl2KpPYm0Wn0/
MTJYK5oKS8sZa6z+SNzf8q+mM4PgsolhqBXM30tKm/ZMHh9FYQDUWRRIeSWm3+qc
DXekP+dPsKCH9O0vxD0pux+bQbMU8kEuUk8UyyLwOx8MTb7Wuz2JRiG/oOew6cJT
FDWbCn+hVWgESUJ4HxoXFg+0ZgRjzTiEMZVuWYSq7gtWdtFN7hHYAXoeYG9ruca5
MT18kex7+GqMBkH0tBPIoWMLJeXEXZhj91+Czm4sS23TzBoRzWO7Ypa78GVZEW9T
jJVhNOuf0d5/8PS+MtCAW5JwXdB+IcQVQAnwC36kDIYwo1Yxq2V9tOEtpJhPg/0T
Je5VM/cLxoiRdd1/3VrCbCphqGnllZoCk5EcSQ7YNJtYbgm5orswarQX/ANHCLb8
K33yGX+v5TGWt1Zz474yA5cC1TE9xvEWOfB/oP0ab1i5hEba/Lk+wT5fO9tw3Ug2
mVqUGa572nJgpj5e6XZM3c42qircBKhIYR+OaXS+sPuvmIEdq8NR+9AgqF8O21kP
nrc/YhOg2qnBun1OszN2qB5RiObc4jNUrxDbBDkigkvvlA51BPC6PU0AlH/lSder
9F+ySEbaQLIuYrH6jeNgDknNIgZnlsOfQDDPxa9Rp2OibrsplV9yAaTC/oiUG/mR
qRQl/BHBZjqaJNh49OwSlJLlB8oUWaXaR/Cm9pQmfUdsHfrQzyzyzqtl0kklTEfM
/PO/3KMm1qcpDNsDV7edzH89vuEbTfk+2OoYuokqledzneIQMNj+QqBilmDYPW7G
zQZ72jKv71XqMu7aXNKoRL8Hg5TDCmsAmEU+LU8Tbb5PRJCeonN2XKOz8YRMzgh1
ahWcWpdQcClu9FTnmwHwjL4blWBS31tDE1KR683C55Z9skOs80+JuCbeXRB/lNS7
IIP3/+B5CroOn35RF67y/umbjE9E0VM2F5BJgG12DkcnWBIUYCjoYUHDUKlX+mmF
nQEMo6Q4M97siNzO80vxJSmx6PJ7z6zz2UP6EaeRMrggeCbeSM7WP/4L35L71YwA
Fod2eynigNvwXIZHHcl8qzo3QKgj/pF97oyxRZnF5V48pwt/fH/7hd2MStAQ2CS4
r5b0W2/vuJGJyH3qT778lZpOvVDlNVpEB6UzTYrWlfIRIX4K3pISTQQ30O5/k8rh
Bp7uwl9vdwHoGcqR1bvw9FbV53paM3t2/zav45o/v8amj/V2My40wf05e8zEmMi0
ETfxMNRSTSszEWnBOFuoyNaoBF76GCeXKKOKHrampm/34tZQNHMxps5xWF39Aw+B
SLsLswhQmC+O6IX3W9694PCTotX6dzwHV6Ex2JVmnvnYHsIU9jt6wf/veBAdZkfm
4SJSC0N2Wh6Z8StYV8uSnQZExclryFaUHju/vlyRLSx3+wzOUoxWwbRu4jbGImJD
V5Qp5l57Ff/fsBIVtFaNcGOwpRCgqTRjhcj6R1VwMkyL2v9ercevqTKskMj3Dzj2
D3ewX8yrpeRM+sBW3jmc3xcEY8bPLJAf+827/4UXucSqhDplY/+QSVvD6ueKZi6C
iNnN2J0z5LSIr6hem0o4Y6Yh/lOIn+WpBjBNooC92Fn9jpc6VH8zOrFsu9rNH0lK
s4VJThfilzIviox00/dlUxQAuiXeMovjtbpjazTCnAWebieJkO8P2FBUazMuEfta
w3g6O7KPkefvwWQ3GRiS7qCiwnh+SIhP35x6AaSWMsxWp6OUZDFp2+OarFe4+j5G
mCSWDtzDqFLmEZzBgt9REixb4Ba8ei/nQJdKxnYRlHLUEVRJx2R97cDjAEHkQ7Gs
j/OWlSyUZbCGWfpMUwaFkFotkGjABclNiBhVVjCxetGmJJWgByDjqxUYqyFFtJA/
QJlZRcoqI0yDzMX9m8RAudTBPfYW7YJDFvE9dIxSrZwD7JoUdIY21WRZLF/1pDk1
G6Jmkdan5UsOPCWsctjBRP0rp+JDd33y23JyeW+h1Xc0juWyS+QDNnyyDAIamta0
QRakTL0+z+RfKHBlocBgv9Ng3jlI6mGUf2z7HxJZv6gIStLvFnc+FYo7NBhsxsyo
ezk7wNY1GIIueLPd7jvi1KGaQqTuNl4qUzS4mKEx2jkV8gCxMeHsPubWRE5cKZez
hRXmHCPe2EkgXlkBp4dMIHEnCUVXvvAY7KF3RusFbU51IUfOjQvgkIPvzNAslJsz
shA3wrtPHOtwIw1Et/M8VKXE5SI31yWLcr6xoOStqvmyMChqn9RLGOnJkey1/0nW
YkWkhOviegTC8blDYeTX7CTorJp5Ji0SgCIw3NqPrTSPheVJIR5ruDjVLwMvXTZw
qF6KjsC7S3yiemnEVDvUw64H/dmnju+9lKRYdF7clUZ1u5k35qz29pPK2dHnzHcm
/HsFnCSde7/omIX3LayAkSCfwBAIRpyFdqQsx4gwhZz5SSVdvhgvuRTy3QHUl91Q
gGBQghyzK8f9Gk0FfR1S8RCyz1ezYr1Zfgku8DgtVShR+8hWzY1HKRiKTzH+v461
q+PRZjJ8Tp1ijneIEbkpin4/65a0MUSqJAIHeD1Shrh00IM3oqTvsYc8aA9C/VAy
Ifk24iErpEGT1SwW7rAWL5+ZmWLHrUKqNbkjZV8wvVNP8Kr6Ue0da3vZBH0rcE8H
pnLEq9VjWReqfRLOy+VXjN7mj7saH1bN6fo/6/I7reW7W1MqbWmqvB8LmCvJKBZv
Xoya5u0kh+V+IvAbNrll5xpFaQNIuxrEB8LfAMyIKOHJ+B9bN/C77MOyKKj6IeHv
/PnarsGs9qGBVpcQheYerv66csDDAqL55ZujSirC+47YNI+/mzoUYebutJ0aCJYd
f26ty0wdFRD3+f417GQWL/Y0p3+VA0pti8YzdQF7sYqsyZGOYwlYxqgnsPblh5UN
XQZoai9ieFRYPqKvNxyVEzB7PSOcZ9HYIoliFY0Y9vYUBwbMSAno1GMJbxBX47Sv
lysIFchAlt0Zy7s05xhRX8x7Mkcx0WOV+xjhoPW5nfRu19Q8UYfeVlFZBjVVK1m6
aDQta1d477n/3Q5YBJCkXoPCCzCYUzECmLrbEnu99Y8j2l1TjZ1/JQmiBJgNyC5L
o0FNX3OO3tOiVuyx3xcSrPiup47Qfs7QMgPeND9Q3r5RGZq/MeXBObznWMQG0FkK
0b56IvS/1ukJNsA6HCJX5GMJ0M/C9DunithD059thvaJwRQTpQZmxAgtTk2l2ISt
AG6MhGxuvYS5Nr5qQTIFpPA3lmk7FfTkWHmXhfQ/kagVWQOFy8vnrg16Hg7QaWnY
DSEc1aZFbLYZCeng/oqwkuxhcQOMepZ/oxsXViWRzLjr9El8hdNC4olCGzwjbCbH
UI1cc1QSgpteH6Y9ln6nZDBoTEkaxGbYPH/gDbFfhBvF0KeANHH0EfpKIBtphiYJ
3rCYIkIdk/+pYEiFLSIKJS0uH0iCnw3tmswb18WoTUa6BWurobaF7F++zAfeVjg9
lBJuMTPoB6rQqtBFVtiP16UYRkMPVPs4Pcn28AEcCB1+9oZADYDlhKloN9+L+ADw
lSIdLEOpR1LWYacvWMSSqPF9bVzSUbqGzfwefIZS/w5qso4XT5h+gRh+mzt+nmCL
JKm1JHaXzpaTZ8MsbHRTEE071PdMz+xrGBQkMdCoVgaLf9hEd7TQs12jijiFikrZ
WwitbF+fL9ZB94OfChsPmMJIlOsi9YOdOie/MKMq7FtxVz0wtecQbPDE+C/GIPwC
8iKoAti5udej+1ZdXYYHstGNMg5aXKFVUoWLvfoDW9fuz0nL/k8WqUBFheuDuzbd
5IvrsbLPfQKiHH9j9jUyl0qz6AhSKN4LjFmau+3B3T9U2tpwoG4ROoCpq12f4oXd
6yfiK0ENhf6l0+xuzzQJ6V8unTfmVppgu/PnFfZrM4p4FYzVkksedQ1JuHN3TXig
bMxtu3zEc2+Sq2QCz4xJoj08aqsHPeETDTH+2L6O/NT9EBqaRYXm4sPpOXqRSbhg
IooMqnMyuNZiGrwgwikgs3aVw2386xWExyzGr22A5/nDcdSu1KiBGlbjofVvbszW
L52PQQroA6uUMWvAqJJp0h0OwuHlFaOVCuEqfawdojYcpQKxAr2VMrFC/y72wdia
Y0Rz+C1nm/s2gtNqzD9G/uAix2KJFJKBoAdskZDfcZdo3BUj5Qun+jgU31ybAiS5
zWeadzmRqxIIvgGEXg08FEAkRU0JVVDA3h6/yyzSLD0JNlwU/hGf1+RR/eIuimAl
YetCFt11zH7Xu/xfE2AhEb0bo+r2JkxVTZCK59nCByuyE/avueCWutymRze0gaDo
k1C422VxUJnONFhVL0Ug3lIgo7RZV22UJe1AOV5Tv4SCazRz1vbGWc7+JN0mVXK8
zhGyIXts/fXP+Ird6qE58zaiXMA4LfeTlhz8pOZuLUR4yKcDZKj0fjtyDnm/YDdW
CjwNFs6pbReJZ1BCKrhH2J2AbsBdKAiptJs01ygiufNc0QmU6e22fkpE/u7Cgtkg
5Y25qu620O5YcHjDGqZ7juoKeBcmf4o/UmuSq7Oqtfm3HvXMJM/3n9RcSc8+mRcv
Da39aSiS+c4b05vPAVaQGwusMhoGnwSpTIVIjMj3oYtOWBGYkNJBF4UiXePZkEhN
7K3uvQ75wopZPP+2K8LILCtTJDR8CmLs9Au1Nv8RzffJ25YohXrWIKRwW6tVlmBo
97IzTCkHA3KxAhEf6XLosNtradxYEUVwg60ZMCCqLQB0lSD7QkYMLen/PAxmXvPd
m2HFnIRUzcyTQ6assJ9/lVgHEy179mVZobEB0n3hVOxIS4LajhsMfHkUZmfKOM5W
kdFVC/EDhRzdEIjRR9pYMByBacob6yIBL83qwFqtMGZfxTg/bEdUTN6EH3+CE2tW
RSYTNigWgtoNjOwoariCbKZjzZ2Z8oX1lFGssv7nf3pI14C8pvUOH6EPwGDyEkFg
Vhu7Zpmas5rxOJKPJyC4eUJUZkcWyIOPLTaBYaAQNsjq775X3AODinuRm3Ot3KHu
sAwK6JuBwO+wj/0sNNlj3OMmtAQ7rNghEKJe9a1AG4dzORyJYKgyWhpPMyTFSrIe
iL3JwxdgWXOsSa0fW8Yi3pdwMK/0whgg8lr1ZqLHq3Rm6ziWdgZH3qehYlRcH+eV
CHEsHtm3p5SE6O6ZU3/OTHHJzWpvoreMeesBM+y0cXcp7iR7BkysFUiDYdepxYkc
Cwn/SFEa+draJolrXvCFOv3z5KJfmfdNw9UVPEqinA9F8/wbbxcbTOdPqpH20w0v
hVKyDFo8SHEYHnBAJbvIwuuBNZu7TARUjLY7KjoEIVK83sNobc4hoEaZpZakqDnx
9zeqrfVgDZBJ0b3nkbDNHsM+UHuUtOgPELgfjyV/Mtpf5gqUQdF9lgxYNh1l3SJc
0hBvverRpFgGRLxjf7ZRjTg/QGNreH2J6GkDMilyGS00r09qn6gJxxHK1yLectbS
3uXsbStcGEF5Xol3ZJS6t2URXicqvLFVpzVHYal+7+5eW5ZPUfF6XVfWueuwf79P
41OujzfaMdTnf0ME0s3aJpO3ovSruklQHcho4IyrzHXeNsUKfAQQYsEgIXG6ZDSD
2qQ4vch7DetOu/7bqOEOdFpFwf+48Pd5Aj7R8QZn4hCzboZgl/pWQId+FoTUOmDZ
2lHqg0NB+XDEUzA91t6YhGh5nqMDADB5XySbiNrQdc5gQQ19i4JBzoaw2oRQJt5j
wrMWH2/nsqXDkKpIPg9JgmZiVJi2T3FvlqE2C6R3GfIk7TD/yEvsZLL8YPkA9Xvs
ofdCdU5YzwWml9FtOSNyiLTC+Lqqlr9AcetapCaNgiwxiIGGMDVCrRt+y7mHetNa
kwmwhzFhjz3Yy+zFCTEazPGtE8PVX/ND8n4UOvOYQrONSwZKn2MB8GOXf2GULwgc
plsWpYP2MkLHc/1EBkJHD1a9yY86UhP2harc8IMFH/n+xh9e71gB5NOJ2uWY0Npw
tLFzdYezh1CMcbbLFmyHUk+ijy/ovP5+Jykd6KwiZHNzXqWUoQzMITmHCkbwvmyL
GT6bCHvCS9cBfuwUrVVVqAFylwxZhS0oj7e6m+01n6Ffg3jBZ7p28WHQIM5Izn+7
ZAaY3Jl88pOqcYfG3dgTciMgFAAqeTdhwT1l0Fieuw52zgUjqjgX7usJ0tYzHZEV
AwPo2iFhvK0t90q3BtOHmK3GfwuMGXeJJGbDt4MM1/DG7a2S8cj+WX88aQZFuEjv
9YUD+jhVxplKCqc7vNlRvyoXNkhfUMtrKbH91qqYSmvSJ1OTsZNJ6HkhW8RKabCv
w4Ig/nzTt9xd5Je+kgWq+qSVPuhnrark51T2UGBOBcoPIpovzFwKVahbh6DtA26T
gwZ97ThkbtQAZIb1RE2rhMSdASH7Pls3JKkHmm6NIAGGaEud8jdZytakFWsy6abL
iHJLKzhoYMCpsZJKimn5Lh9vZwpBaTznBHUm9UuWzdpjs6gYtpOuyQK8RcuAteTS
+NdOeNoKBRtYqI8XOBFrI0MulUN0m5NbV7D29mR82Zz1GJ4okmNUcqeDOAQYErbo
0hfMPlE33vzWw2jQVPP4TzfsxyVsgID9Z1ZGq22SYsV5ZE5sfjVpYN4xdM2hR4Nc
oXXh+UI6En9Wg5GdY4v1owCqvkXknubgS9Y+Fi2AS78wR30ZOOqXijK53QE4jKcn
h1TLCzrs+Mvh/edZarKNnNnP2NIFbOhikiB/Ehv5EnfmvZpwL3luCilsgFpRRzKW
Yzk1c4LCpEv4YZkVlcrXgx4DlnbQSdEAZA3zNbmJPFelOE76paJFHGYKQlYNyOoR
Zdix1vIdyqDE++KFsVxuRNjNq3PizITKvw0KZEcSrVqBuSMmwaRqxLBWaW7G9cok
dVqMHI7DSgjcIwKrONYSTrh67x6WAw+61G9EAUyJiuiPg5UJc3Q6worlH5e+uKc0
+3JnI4psrFRyc9oHsBv4y5V1YZY7NQGTAvbnwy8pqiRG9rkbSjyU8NexFzgdWyi1
cJqttRIAAeKEtV8mqVguIhs88PdIrGx4ZENMgC+7qsCbIj/SYe1Mwu+PnQ/T4ZtM
5p2FgAwQRmWqYwL0Eo4qfLPDB1LfvSP7k29jtHKDeCCo63VWMPNJG2ttybJ11pfv
d+zpoEEpFvjKqDcXIdgK6JhQh9CXonSuW50uQBDnr+6h6YSvT53HN52tZFC+ExkC
JKYUBj8qtzTy08djXz09nq3iqc3mVglPaNC+nTmBrbQ+m4UgX0ApGjxz4ctp2Sf+
8feQJwJbT/seKFmy/CFxm7Sv0KS3kmIyif/7spNJ+wFqBXwQYpXBH0DCc186YOaH
iwNzfIyT0juavvo6HTKcmDXOxZbbSaIUny5fkjKAtGOA48hjEdlg2W1EeJs1BzGo
vIqankOdXiEMkG/wHgojqL7puG7Q4l7KLKkw19u2ujwfgY5F+57OHNNGS8v0dUqg
/10Z0QW2n81WzOQpMkmc+epkHD72Shm9yCrTODLc0opC9d62l5uW5ocDG5s4dCZe
vh36aJ1hlyGq691bBYWs0n4kGlsTMsA6GDftZLEPqENb3PM7E8fuvlJ+cD5XuJf6
ZfQ3K5VegSrh8PEQIGfk0dcaMnKWI+DUK6dPfZDob5qshYKSZ9sS0LnuOzPEeID9
1rRubj9Q+oYwmYr1WYP1CRwjEutgnxrmfPGVqqVzvK2+aW4eIHc2pseokbBvnyMc
VLIBPrrh/03PAZUiPOHHry/AjhhNtqPpTUrKvJZEpEauUM8yCdcKd/DSPGwQBK0Z
/jBP8qgqbe7XV8HP6/rfOhNiTSo7YXv7lHqnBY/XbKPr5ZybTZTwPoMuX6yjvKXn
AvEOrI4ygIwEVSBQj7b7QJhDYztjL4RM0jNuN4cQE7mMvOJMVWkcmhQHddZHiWgx
Df+pMNVcTcMF1/xW1F1ujNsFnsrbodcNXJh8cL7DJcSm33R0GxsJIz+3Z1ZJ+Q6T
RrCFfQmh6S9xJY2Od19oG+xltQoe2DQ2tkQa3RLUr4PSFlxXWVKcvLiVmTxTsvBp
7hRjTZYVe1I3KFYpZYZgL+xerW/W3+gj5kjQ3WLUOeg8zzxbLxQw0FMLLcrHXJC1
ANjGAqM7mkqkYaqlahCGCjNUWkw4ONSeU8/CxFK3VGW9iEV65XPeiYR/CPSGe1wD
m18Husxo0agIQpb2EW1bBmTClvwy5Kh0wPdWSuNH3R3oV2MbMf33/wMc0WnaXbz0
32ca0dUOpIA933zvPVbQYYIPfXQ+5QyqEtlVGt7aljXpmIQXu7FcdEgJNZ3WfYPj
vhVcwWl2Hnqkk2x+R/vH6eYFKW3/KBjwh5D3qD9/ZQKDKxvg1ZTyHE4imHnqJro7
lGCkNN6vrRmN4f4pFiFoovtv1c2PLyLD3SdokRQhzz1sCJ3hKcRRsypJVeXl2oyH
JFo/ts6xiL3KdwCnpG5mjchayS3MMOpE3QaOB8VjnuTnEP2yG+CEp/rKGuUq9cWZ
vtcAxxCTNYe7cxcE/rXORW9KqvRWvdOhJvjso0qq6RUNYhGCyPcUsv0+daB8o4PX
qtkbU/SIQofrLvumftHXf1soiY+iq1XeTMQh6BZ8YVhpzMUrIrCuXdwBp0bmEN5w
3THl23M186pMuHBu27imuurWB8uJjtYvGadfW+BkchyNNJBZNrE8O1vCtxx0b397
hTMyLGcLOFjedivHwlBKstL9FD2sr9rqzysA0iv9EYdsmvt+wVSacDsjuHU0qudk
BRKyPKez9fZvsxi2vO/cjTMqkeyP9Hf0ZzAtWfxq8BPveRWxwOkGBa+lNOHs8TzC
KTPYfZRjN2SIxscAAEiS6EThUF+ZqoNWKvYE1MZnLiSEhGQSCa6u4wo2fs6AHjvr
oVNdq0FjCiH8WQgaNN2FqIzUAFK0kM5fb3+dIyJp5gZj6Zw+sKzXOEkrkO1S1+CC
+NHhKJLiY2DX+b1E/LxARHHfYerG79cnkAal9R9/y2OAvmcisn+xJ96S71Hxzxws
DcB0Y3Zm7eFczou175jGg7ecvY8UW83zBay9XiwPisYnwISkSksaCOkOlhkw7d1x
QZ6t0t5qoEI0lRM5swCRLRkkQtMNEr500Z6Bkdzc9tt+Zf6YtNVg/Xid9A75RLPP
b00Ekh0NYzp54iEapf39cyasdVQwKHKexb9xmuPAFJcSV4yDFlxJmfr/mrBwlqoY
n19duJBEgogMHce4/Vcf8Sll4Ut9myQV4Ymn9xESPZSr1VJRZ6iZ8hpulSblxdmu
lbb2MaIAhDU2/mK3Oh7iSCGeQMYsTayGqoteD4Tv8sp+0LanBbbXfnQ96ZOPA6HH
QLmoAl0hO+Y6CwiQ/1lcg+5i4R6jTOkqHff3e1r6gFdu42CCeRzlp09X926HMzwN
iMRQ6dJTzJYHI+7Ym5XF8xdRCOmkrDnG42EJ05io9faWhzG9SFadULIKzDocgbt7
TguqGG+6Bv9sTwJxOYhOpQL9KEVCtGvSwOFCtqpkL815DgPACvvKUf1mB/6OqMiV
m1FfQ+Xup2PSW4yZxV/C6G89GqTA2vnjCvb8f982VNbRKPdCNW7zurkP5OtPQlDg
EYFVQN9jCyKTgnwVuq7hzJhZsCRYe6p8sRabr/JXhcLsAwDSGaYp3zpqUcGmd3eb
nS9PtyDqDTFQGny3qVV/w/WnO1c2AoARBSe/0qZ/4O53DijGrK7yjubyLa7DqTlQ
IXddUsVzD8+r/jxgGdDgr3e4pwj3AN0FNFlNXx5BMHIwBBC9qZ9eUO8ANB7sDB41
DQixlg2Gj6/Lyq/SrJtg9Oyf78fnBp+iTqGFewVTH8JpXZVxN+kU1Pp1IL6wswHr
xIwcCFMdYDMntP5z2iq/qJrJQRVKuuUhR6ae5zOECQ95PKtajDnhhLSC6BMQqE3P
xZYhMx2V7QnZAaGz7+i4R6wX8RJ0Y9osVM58uZqm2MoGPom3w9HOCVo3kZpxBMNX
MeNkeIeNvqAyvpbT+Mgxthpl/G4IyPPTCNREmzfoJfRJJ6zoaHBOKaPJoLI8MU+2
ettBTD6hH5NWaEiecYYkKESNp2m14Xo2SqGbvSKPFMibAY/vApjZ/pDgPH1yTiYa
g2gfCLGpOlgYrAJLGRdsa8REFEVp5udpxpyJxVgeN/Ucb3tQsElSsDbj/q3+IR3F
YX1kGPUIXO1e4Rxdan7EmsZm0hFu0DQas/ZTCY2yJE9vcQcq6ovWxMt+Pm/l+SOC
EC+btEUQXxTSla7t2WR8bl6Y/EIdBAp+P7Sh8AHqpkFCAbgm7r+iAVIoNl439xv7
p3DZATwpU/ENwCkE8a0PySR3VfWH29nzQcxoMIno1e+g3f02/3JixXi2zI+Qh/BU
xPejM0hv2cgt6B+nLbN+WBPr0IycYDZou3eCopOaHT5yfVMJ08ZMQOJHgdBdWwH1
NAg7M7XAxxujAGEUDD9XRHiue5aochpGNPK+Bg8eOmZsvjhgdM74kfLdpkvVQy/f
09QHzv22JYtdAnpiW/cgz5I6jYZ3vkFMM7z+hVCNVKxvvkekKPK2hU4pZQKbveH8
QZEyDhgyZH7RKbUENEyIkZkZJq5J3NJfU61iJ2Yfu/0rmzZmND6flzAedfI3gFYW
n42KR52H3tS0yhZugSUtlE4CxBNhtHEg4+yMm0pNlvBJSEgUloYHpLIv7dad2yMh
RSSFuMF8tQ2AI/GiQlwlfUVBDDeRu4aAi9ypLdRS8BJjBV8IeE+BDMO4xL7hg+oO
Rp8spxTAsDO5KvD9OcSJPfbj3dhm4Zwk4uyHmqULrYBRthMEQCe7XUo55BWXuah4
tQNWtostuUcdJJ7tgKOOcAWk3szJ3ayzPBX+sGQx4Y0Q2OOQEWmEo9oYQW46yWOf
IeuNBwKKZzSPHR7EP0bkOxCjEPx0S36gwo4b8ZWt/fsuhzhJdyrr09naE1ysAniE
ACLc4RltYpyuA3zYVDQPml69e5BSjRqY7F9uxuSO4tPhVzqKXYsmKcZLRjNKv/6t
6HvtLCwejh9CdfpnAjLhLGvX2UxH8VN7nBZiIVaAjf1fDXzt5elJBdvLQhclSvJs
aNgVRM/DRQ9kKviSijIbFSn9dN4DYyOw9vSuKcJmVRT10q6Z1kQ9p7C2vN1kqkMm
5MRbq/vX9R6gSWhee3wPsQbF9lLtkxKeMmKUnw0oyW1s3KUI7H9Qgxd2f5V4Gto1
mGsjM9XeyJP2dUPCsTTL5vBhiABEHqUPCTlwLdoHqMhcmc8Fjq+4rUZ9g8E4f9zN
wNf4h9yQLmZj6Jpls/W0WPWsx7i74pT1Bnl9b8xC1TsmZmpqzhyovWlU2i0GZn3j
85jIHlWaj2hnhQX/Sr7i0F52HjUzVEW6ln/KtBmAHqKo2alMzPjwmG93eEegQT5r
xsCZOsxWAv6D9l6DyX77Qn3XzX4qpnz5IMn8ZREQPFyJLjBVYBAy7HOdfksVAUlN
TzRvhpWIeql0aBofng/7s0FbhRWnZtgtN0T1dGJvHD7jv8Hdc866X+TjRfqmjnrT
9OxvS0A9ySDLe7/E4A0N6OSxgNyujon2ZgJNeq2XN5To8Txuapaby5Eefux9NgEC
LF2Q76JPFjiDqLPCYX7xsY3gyOd1JC4i1lxib2pwzmBBTJoOpVgLMHmNVxV/+P+l
Z+yQbddSymS5Aezks4T9E6qq/QT7fOgd4t6fXevShaPTu4ltlf5tKhok1QoThyGr
TcMvnEKJjRxxwUXlqLxOKT81G4QpyA7b57WFC9dGPFLvueEEVBtdpYziREzfx27+
HbXzm+E11yRoiDJF1aA7Z2AALyEem73uJBJtClbBJaSTuS/Wemh8c7GxqaDxfj+U
+Szqy/FfKkn30++sWZojahHjctZmDTybRwEbtLveD/hy+oIAh+yHeqcZdvd039wh
FEQOMeY3aO7uJjPPTdJ3qf4iyJgQrff1vpnc5+meO805w5tXlw6VFOEN34QpCERn
Bnk7BM3MseLBZe5j+6lxhDtL/8oX5GbHX83gi3IgQvI/FDzE7+Ee22H19SOE4opF
aDyYe8amdBW+QF0Ui9pi4Qq3LF5+kxSaoLLTpqddSsb5XMgHhy9nYBAL0/7/O3Bs
TlqOwnN5jnt6JiketxxXnEQMWVsU+WTtowote8RqtSK9kOEvVNwW0aFxwSp+ODMS
ZKJBAWq3VTv+R+EZBW1zg6grX0178QNt5bWPH3sRhIMnZFxrJS0LfDSxl6BSKbOA
i3Z7kR6hXlU8/QnkwN0VYiK1OeXap3LaikvI5+53kuaBJeDnGu5oQxnkkL8903FO
mE2VnnERamDB9RA8aIZdQ48vfnBJ41wAP5pWkYYXK8i4IbAIu+lA91GDy0UYlGeh
Fxn6D7DfJwo4l10+kEuO5HiAyaSNJT1lGO38AABjQIRoA+LfMhVYrqCEGiC5PmAA
hgsm49kCrS8MMp5t6hfmcSagp8Si1odLS3pZ933E1Cx2zyJ0BPUEf0lDafsV/+Bl
3ctZeO+T1AqO7bX2y2ZSaCZMzWQfhWOy7bL20fpHlf6PRKQt0yXHIsopkqzLkFBJ
FebLVXeOu77Q5sDoNm85El9+/+Jv92ZvrJ73UJ+KNY3HZPEjeMcTsRnvRUpx9baw
BovhZPKmixDibd3drA2MbHzLmlrKONWu65VqXzaN56Kf+6hAK7w/GlPFMhyh7Xs/
y+/HSkivQMj3nlpATllE1XfJib8Gal0s/KgavOLewksEmIFbYM9SHKUR3njQ/SA/
9/QHjT735ur/yuYGxYHzqRTH2k2+dEPtpoXtRXgUtby2Tcuq3KoJfe6nURxr+g21
DpxdB3obe0BPNMnuq4oGVgsCel4hjXDqbKmsRwXeKrNMHn7m4pSyGCOgf3jRHgAa
didxeINhhdlUAUb7b0pspzaDB0+8aSzMkMvgbD1IYsRrejVidVq4/LptuBH2TSuW
wC5q2kVuRMYET0plBRHxa2eW3a3woy4cbpXSgdmu81feueTvQBnkw2GEpD1Ivwf0
7gxXLECOKMcJemC8srrG13mBmpzJUHbBCcQEmgqtyGxMbPchhyl6No6jkdOthaA4
CkxCqS7DSzBaBFELfMncU+AauPd01W6i1gy+t/6kZqzmnprDuS6nYwEFE0RNTh4I
z6qqeGfOldaHH8wacEBsIksnPb28yu0yGMe7AGxkcr7D6s0uo/0IPxkestjyEP/v
qmndZyWYItODEaGXjxMHlPzZn2LYHBmtpfariJ6Xc1QUFs/M1XVf3pIHkkYG8UHn
NzH2ije7BOlA9Sk8AfxTHgo7T9+bcstVtnS3y5mX0OzieLkiLfDJIQyWImLN+b3V
APzVspQuTQgblKMhq1SJaycv4qCBKhaVijunQWmXqCLQcdYP35iKREfJexHqjx4N
DhA5NqIsXbyZudsYFVVrlWqBtI0fBuhbpyS7mOgkFb546kOvuWmFu2S1nNvqIuAP
ZIwhtf/AnTXYitLYgBPmLPsg7tKDCJFkxkzVAjEZWSRLbgYrzMd8Q3URk39Te/Ze
xsYbYwroHCVw/p6U+P2nMwpw1H552f7E8TP7XEBGk3b8d6R4wgB0ij0AV32q7Uwz
HSzo6iJGetqmvKrcKUIqH7ISFziJUwpB4hzrk23yYqL/FnnVwUc9NTSnUKHSjCM8
2az56C5ulHm3dtGuFEgg42gw2Mp2fJyF7RuwfpGoNMx7aRAZt73INrP+0PuJy6CE
ersSnbS+ztQ8dRb9NwYuHalHPHTKKjcn4SMh9O9aiemQTwReieVBE+qr+RtONby/
N/dpnnknoOAullqw+vLowbpzvLn+H0Bu+LQTHEaMPowi8GyBaKcbqBvjuUFSVAlh
pPVFnimDJzEO2/13REM6Q6Hv2H4jJ7BUCMvf0Xs7oEx3nw0FerVgB09vbyL+Pzef
0MeRG94fSplVf3zf5SnN4XVocZO/Znm2JzG+WPcM5rEkZuUucgiXXjqZRW/0DSIY
8QuQXWF0tZDEp4X1rVck0AUPB6wfjVaA4q30KMfs/TxYf7OvDnKuCD5li+lLyZWv
kBV7VNCURpj3xhfDN0VzbGBSjT1KP96hg+f9ZoOS3v8kahVQCMLCOzuP4UMowk4T
85jaNCJGvBGJw54AP1piak04mD5s9kzlzyNlxeSPcMFmEPzYeRpq4sGk6Jk1K+ku
i8AwM0SWTT8otq1ynQu0+MAd3iLrCcyIjaGpy5ifhSq/QQEo8zYrZx3i5H4MymeF
ejrJa/oBOXMI4ofBTVyVeUrievAVCYt9kkpeq63U8UOhbY9g0D5gCF4nBoGDAHDD
B7NXLon+xBcTq6xEsiI/4PnuE5WtMUZPuH21Ev5hWWRlU3Y9JRTXBjWnsZ2El7xD
pjXCsypEHjMIa/AFdkkLhoq3Jd7S0oG9KbItzsAI/bflpmHcEE9x4qiW4RZVVvAT
EFdSEhqNDok84wAwAoljMJgpEWTOmwZ3OTZPbNvpTMKJTGomI6ERIMSoDAUyJA/U
Ir3ojaSg7ZihYv2KUCbSX7G/aqbueDpf9mdhq0+YDRwrQSHugkLlRpIt0hkj0q5J
CDC5i5XKsQ7WG+dEJcKQ41ba0dot8jQ3Te3TXGpFVg9qlq5RFVm9xxjveW/W9SoQ
2NdE2b7VlqVOkMW4gIVMyxTC1oNViHFEgVBgVxrpHwj28wt5eAG/PLp9SV9kfSqG
g9Ki6BRAkwCbtxCAhxgyiFNSSChxgH0Ylp1l/zY0PcnmhxeUR4p1UoBa2xQXm0W8
bk7jHgaWtrGAOfcCqmMNYzOGZRQPyngynEA6dVMfrjX2toUE6PEHz4PPKLWU3bPt
2fNAP/3g7lPjjY8IdSQAIX1YpPaOCLpyzf4yg1p9yPJw1OpAg3bLqUljG9imOOGF
8SGf3zXP7Bm8YJX3tTd6TcAtB/wgHbPaxfy+0kcmQKVviYhw5IGVg3vggXJYvIME
mZyVZI8o7dtjrWHKCwgr9ZhnAoizkyDrhg+KioudtDwsGxzeDVi/4Kq3OqI7wjki
jpzlMDhEgDp8/M5MBQXGoOPf2ppWCVMMNPJyklts210v0ibKjawiWpsxsBaZPKYr
hrr2jaZ7xtYx3c4upCt/qcqfAIcRC4VU3m3GOWoTfovn2te+z4V4rTJc10QMw5eF
yb0CNzTbZOxS0wTS9HK9ICAwrcGp5dzJiVO/170gz5w3A/eyOShuW+VCr3fAltzQ
9t6c1SaH/aWFThNPGPXESMxUHp+HP1fX0v3IgK9jGvx0zjlKH3sj2RniGIO7FOa6
cetpEZLniAXAfdjgm3Hz2APwXCiD6eIrRg4W3D+wG6WwmVPS/jkc+Tu3iyUBR6ho
0bpuPsQf0QFByFqLttIOIJO7H4O+wcfx8zsVWN6NHp+aDD3Zq/YpIXR4ULCGkpcE
qZDJ+CZ3T1qd4764izVatfKLZoL56aoiXjFu8ZN2zVBL9mbA+3DmZFEEgEKwCP/F
qOJgK9JL3afHQQlTTE7BC9yjuS9Yks8BXjtoXyNPeOE+hWoJqx+Db7Nyio/bdynW
lGbd5U+i+EwDgXf3bDDxhaNyDVv4cUPBD/t6GJYfZQeawMkl1IWMks9UHG4xrWhh
eTFBE/qwea0fAknqkX8/StVWzabPleuvBYN3vwWEbQZnCfYMr5wdC/j3UHEK1n3W
UiryVeq5WArmiVygtQ7T0ND+IJOY8z5YeLj8HUMCMpBo2bT2NHIPnxP0rr0XnFq/
As0TMpA9IpxJHkyCyaX5pae7pA7qiybsiJ0V2kPaXJdpaHuM2sMXFgXa5/KnjhpW
2xnEm4IGoXd8eSw8Touz8xzzLhx7ICUGsDUN4R0VyZaTtatkV6XAgZU8xbfSYFZX
vo4Li/QcaWIUB7bN5VuYEHpBaR7VkSCAeyM07gJg/lahv58t4P2FfNH7YoKDnmuk
fJ4h67/O2pHiduiK3MmWaKKOIKWSIHnr7oSax2tFOtsBdeekarVosfCxagBwN5bO
YqMcmjjbyvhlBKuRZo/XztJ9EGtV7bYz8bgDd9YUguT4N0D5S9uQTUH8WNZq7lyG
6Sh74TTexRC2+Ze8T6EREYS6/aLbekdh8n+RLdqUiWPBqo5zYaZEBH96v+NDYP0J
8b3LrHQVABR6s/EWHtPuN04T3kk++kt1x8WRDexDcbeijImFS2/S0mXEimwAzsG7
Aj1yjyNN7alAO8gkm4SnVdqLM163gsKyXKUd0b0FpUmLpAeFshTHStV3JJ6iJ/v5
4WWzNlghKSdq94mUoTLOmMMUCFIwpQS10wfY0pHQ7Z9qQR1jnKxLgICfXE7b+jko
M1MIJZHOzz71R4EJ0pt6+u4EdvIMqCKyZ5ELLS1+dtPZLW4wRAMEyWmnbiPHsMLR
e8zT2M7UbedaAsE8CyN6NpblJIKEx43Nc4Ueyh0WxyW6AUjvEQ+AGPyeh18my/CN
FwotQ+FLM5IuEzWiyw93TDS8FpQ5QRChm6hhKPcwFXk+aSrQuav2h1XGFgoFPX9P
ylZ/X9A1vIXJgC5kDJqbZCF8Go4+XJU7figluivmhHnw/rtm63/4iBePIIcUIbkI
K4Bqbc+uVupuuewp8ZYL6WvVyEiNf0sjwNORZjw28zY5rombaQhlGxujWGwPwG3Y
tKNmRpj5VRhfKq1WIgjQFHO4UOUtAGULiqCGvP5DSC6OON5X0+UeLcALc+2Tf2FQ
tmpun955ElolojUu03DzZX8tfkx2V11vf4fA51vZiC/msRzvC2gzCTIZwmDyaU4k
Ps/RQv9CwRI5kWBtAf5t6PxgGNbFfHlYkhz0gfMDgAFFFaulprO1A59auuv7SCKo
1zWvSB8yYEO735ozN4Go06uQm9oQpL5FQuPjRhWiIHRW+hUP8v0mDkP4FwNLXIJZ
mzAg+r+LIclbEVoJ6DdLjBcp05hrdq2cQ/iUZwt4XU9x+0RkiAIZFWAY3clf02uw
pBrirvYgsguPKmCF9FmzTQjCb2uYOun/mSUmJxgrWXq4VII6mmve1vnK6lT12QPK
8T/aNGe1Cl2A3en7rmaklYM5Rao5SS5j29SDBSSkKZcPXbpXO/pLPoXgTZOWSxW+
LpTJFWTSJP7K+89arEr6LoyIuE7d+Mfs55HVHNl6HDeaAr8SET3fQ9on/NNPU6aN
rmR0qKooETceU0uI2FnIjtw1Xz5uJTHqGCAOZL3J3uuTcYSKTtP+Uxo9pCy1K178
NYauCn1jvBjGgisbCuNCIwVeG1Bva9ke4Q2XL2ly7nzg7J8GyPTCN61Fsgdz22gU
vVhft23UwWd5jkDx9huZQm/i95wJGq4Yls6z2j6gIMmjq5aPjKZIyCj/YK0RVU6M
Z7oWbYBgKCd30qHLGRPJkCaVCyMxPsHoPL8DnV5geyp/jagUQov8EWu5QpAlHu04
t0CAPuCLFlHdHc7qn/vHmIS+8HgHAEpo4FkwCpl+wRcgrRiiGKqgG04YnPPgCeD/
VMAQftIvLHxRDaQoVrphw+ZysF37GX1OBIJ2Ae60nIoYxoW36XlV7ylKvfd1fjgx
ALZ9Vzyp+CMF07pEc3EUDTsrH99GLZYEMgoGIeLi1jSiSnYl91Zy07VogpfT2h6j
Owl6PctsIk1GL9VUKhV46QhOWf8zKuE6FN2cqO5LcQQ+vIiqwskSuoNs+z0MFVzq
jq91nK6P4DUSCOxG2UsckpF9FSyLLYLoiVFCV1XwRP/bWgnWC0oB2Vsg9F6jCx88
ZYrZu3w+SvoMDIAq/A2+FLRCvb4+5B1Pl8h9td7ccHGvWJrKFo7pqk2GHQ7RJD6X
9wmtCXXdiSBp3mHCeAD8K556Pg+emq5EcmWheFHn/i3jY/lnmU0jnJNi4mSXSZ3H
zpQ7pOFIbyfMr9eb1xW0Sag6Wa/hQDagsCP6Bzoq01OfQgFYVMoDtrYBZ0l5Yyju
x+pKGQBexYPO34vGb/sJSdhVqHgsyADolXafQfAWQXsVhcfIDcfsi+wWvIQ0+mBN
Skt31ftlDMKW1xNMcN5+vYnz9ZUkpgidGIHvmJjBqXHFpTufGDgBZd9uslo/Mtah
LZUArFbsUGx+iVp4PmNBjnesUHXW+7ybb1qL4bvoBjiyH2dgsFr6fA8TE7R/lrUk
MOxjFFSvjWMwYVytcZWWXwx8HKcOc8lTXl7G8KFf2YoHrW9SgUmF21RgIt8yiSp4
0hyFquVPcQO1ThqPscgVIAoNRQmNepOoOiqsk1eSxYWFXBZr/vfVE3P7d6CsPpdZ
h28wKGt8Ss7F2Q9JewEqzIAnAY3/EuLN1l+KfrtuYALkGB6Y5CMxiQKEWoYP0B5D
VV8wvB4dfF9wwpo6c6Zj5UJ2NB8aGb09qrXEC5954dtvCQiF3VGOtvlOauTfy/uQ
ylpihm+GhBTwxN/jiIrQMYeEHeKvyAP+AjmMQknJ+iQx9oMGSI2ID1NvCOqiAQXH
x5u2JCAYtl7fO3ynghrtgAdNYHYKY59FuaJQKrYQ9Z2grPCxsVZhGBYhUn4OkBhL
eJx0B9a1+wzjmUIB3cc8MLZz0cl3/9IFUTUzpWml3AURERWHq4NfdRR7Mx3JSHRi
APiBnKKgMmIXsWeYwUHLCn/qDwzGxSfOPjuI7A5zLDkPgj2kD3TTZgGK7klLZqrH
JOIZ70MyZ86hXE7PtLbR15ic6aAMoSebXKyRvoxHJlePG+mifWEnAxdIVGFwXH10
AV+GLBV3XQXUV6wYR5ghV/PHqJJtPHLvToP5fHgJiCA6D5MLzsKfHjwp5+F7wrD6
arpYb5SqxWjT9dI9uhHVRdrFTz+YToqZrBTAW+vqGVkiNzSsXc3klKgct4lhmF9e
VguuPNU3wdWvoCIqHHknFkJ0OFC7WccW1xvcknJnzpibe9ZALp+fPBIJf7+iOGm7
W8skRdG/9f9bQJ67V4gEwCtddORe8E9uNnhItNJOlOCQFUQVcp4wVUrv4Inq0QNv
dyqYrpqSBnI5p363iqR2u8P0gbDd9yRuZBseX1fy+0vfE/ExFnZJQ5+Hrqf83FXX
0SooT94+g8/aVHMyOo44PL4LRGw3nyM3mXHmtmM5Yh77cpsyszIjW0NiADjHaS4k
R4u2qKkWJPYbXREuASSE5gqxv+YuggwxAufNYG/a/S2h8hK6Ey3sOALrczwRvNTy
5okyROmia2MZS44xB8NqxL0mV8heHwxqQlc8p3oWDRb5ZzhpR22UccRMx/6qoYME
jhnH7WSBRLVcQXyUkEPy3Abf/KjVLnW/8bNyGeN3tFh5AFWfWsrdh6qbPMLjp5Lh
sZc91/qiLiV7NpkBHLNANcO741ICZtwXbwdo1laeOO3w/P1ae6PUn7ZK1PFe/J8Q
hLtfOdBCCNtgx5lZEuMWrPi0toobGpT+knd7Z/ehZv/bYdwk4PYutqW1KoBKhlUl
U6gOTvGKMuqXp8WyRaraqSedMSEOQ0ATMby+h1AIzpglXCGdQBqwAZ47asyQAvK+
OL9X4Yj4Qn+EwG17LbNl8DLFuI7NKmb/BENOfjH/v5CvxRjB1IGM276367R+yIzk
dbQPtV34ws2QxlwAvVUXIef0blzmH/YxGDeEFKPE6odLohwS2NJb0Q7ZQ2xTYTdy
l1MiXG7L+63YmtXozKJgqx6/8cF59UfJDHlm34+rMt3WGVjj07j2uPwWBMamWJEl
RM4KGcwGExBujKPAQ7eUBJVh59th+R+n6x3ZcgW5Brzkq9okvXYOc3p9W53L9XLt
HeF7ho4jCpimYx2EGYyJUU12d12qiwyvk6sMwXq0xZGCfQDxmJgPosFkDp1a+T7o
ULvwshbFdfl1BBO2mYMTvtqV16xJLuUWkg95zDd1+Ux5Hwrw24HYU9B1aCKQVCrx
lWobhznvesbSJIXPijm04PTBEz4D7Uvb3JZDoiUG58ShMxNdL6oeQmpjDs5SBj0e
Jh5bp6VNI5H9myh/rMarYrKXXuNk7e5pSLZ7uE8FUFqbJZm2SLaVUJMJbfdQDTab
/oDajapp87jFW9A+sopnUoFsBGnEiP1GT8Duztx8LrTf16tmdPKAJK9O7MtNie4E
M0CCKjKzdK/xHyW3d+t4oh5ZsZ1DRZt6ooV1Dd8qS7rI19h49mjTRFJcRwiE6Pj3
LeVDYqy2W527vr92WWSI4jpZt08yq4iB7lpd3KwNpKuQlx7jNziABHHX4H+CQS6u
eOZIt1L6Xs6PZZ1WqXPradPA2/ayq6LZ4byPp6me4SZx5qUhWw244wwjeNvvfOzS
iF8rQlUbvXDeGMAmrT8Dmj48XOQ3QwujOhVUTzUI86d9bEhYRek0j8cdhD7X1EuP
ykLgn3tbudD3VRuJoTBMVi2jZqDtkXoRWQ1F6zZWQ0+Olw5Y5Z0LjQCyKP2nNY6b
/MnjsZG7m1oJO5w4QWBQWiUmxNgZZ4/rAh8FVDwXPSY5xkX78KfpdfttYteTVaxI
Of2xO6x/Eyev4sLpOFnC3BYHL45CS1SFAZ9aFXsXULmlNpNGkDPjKl26bVlueNU3
RNaHJZU3bVFpJPZ+Sw/c2mFww/fSe2yFBJr+r+Q4qJ/ngBzZmMv491VDBTH5LU4o
CANZqk9zCFXO8yiy2pJ12dEt3wKZd9x9Uaih8zSGbi72pMfPRoauoWLwI40nmsQf
PKQCRxuFBx39UowIaCk9YJ5eBxCcA9V8DZbt+YJbu929D4qYT+G+SrGcAcenp5iC
/wjj8eyIOCmMbL3NVDVOjVZuFo/op8wvnLvTTZwkPW1dMlcEFDEbq/Xw1y4paPQd
nnq1pOvJ9iNbpZPWppltFx/ssEQpsb+L+XbFOcrJCQcVcmfctvSXdRwA0F9CD+zK
VjHOqFIKanNCM73yWMUtnnEVOtNxFgjFaMKaCDUS+NCVD1PsLptMSyc/RFHM7Q7L
SngkLE3SVUoK807udTm0uwR0kKAVnDCSYmsJEjCR49t4ik4fPNNvpK84KUwDeadi
rwodzefHG0BZPwKQcVVqXnLq8XL9EkPFRighoc4CyVvNCE8/V1RrbcEw+m0qA+Z/
tO2EVmGnfDBhkkusqujBbr02pVVei55B5I4FidKaq/R2ohGF2XB5LhMgFS2/S0GR
ZaxotEdKo0beS4cJ1vZsgmmH7qdK/WLPhg7Um43tqA0oFgTZzOQLxueqdwmFWPo8
3d6oFF5qzNV268OvlEsCtJ+ODD6g4dIHzna3o4IPYDhcHCbE+eIqpUEzJtd7v9If
fhCwipoxQU7pISmPCyWstxDrW6ymB9XRrLIcPQTGcnlpAMH+INgViLtRkrz4FE/F
1l+F1asMcVXyD5xvbv4btYzZjZJGcxup4Mi5Bh3ojgq7qE9msBPBXDvcs/5QOHpc
KH3LXUhgL5x4XU08Ig0IukHsg5nOCgipmqb82AEDvsvu/ZDc1KIbQusoUP0/8Mhs
vDB+ABClxvW8Oom2fAGfnr6cM05zFWR5+m9bLAPX/HB+hwvWw/CHTRux+aiOFQcO
Idrq3p2VR7XkgyGbhGn1VAGy4Xc0DTfnwZqcnwU5/ijMX97CPh4qNHN/jwSu9ofx
2wCSbv+nRXmiilf1cGf5nMs/M8MoOPk3bXSqVKPwjLK7S1aL357r0Q80vl0zAUtO
TX0tQO0iI5i/w5FgTAtmyzZRyS/BCY4dhr1ZBLYu1AnX3GZ3KEabZwaB2yLReqgg
nQtX1X5TxyhCqO64sGo5+al2l9npfn3v+nacAmX4264BaZm43t09M9pNbglsFHZ+
HFZLpwCGVWWlgSvtU+T2wrudHxy56TSgaX/mQDczu31MR1Rcur9Vg+98uAhMhfLn
1HLO6WxYv2ju4pXpkTXxceDWdXSiZ+geIWq2fLuAw4rZivWwx807nmZI6kOy/Mbh
KsoW0opvwnRwd+TZMjLHK+PuFU/r7vVq4XNhQCpGe1UTL8PK3VOlmAt6a99Pnfmm
/K4ob5gFzkciedFfTf69jgY2zeQzQFA7d1E6Myttycs4frN2e41gs7Q23mGHahmg
/tlPQesPTZus5UAfDyolI/rlbutZlve9A1uvzrzyKGWfKHxC36oRWV4JYmeod/f8
VNLlJ+gZ2aDxtzuyPgh7745cjKE2RVKUJ86XIcFu+oqvLHAcMXx5fu89elphoaHU
VuzUGR3fR1493HcHwzuzvFeByOarWahzn2AsubB0WoOzaq2bVU3+j/JitiQvio5A
I4rnafw1zzKCMDjiJBWcp6R/SgNwbKGKYtMK0shjBR7hNnFwFsvSE4Ji2hN2g7AD
trjBzTRlwyVCp/6FAMOHvKw6lzH7Btz7ncZcY1CrBcyFs2GUXoHqr1usx/RwD4os
y7HKX8ugqoyhZlCwXAolFkBXn01ksjxUvH3qHrZRNW3m5i35hdbcTsGGjEaLHMB/
PDMy4aCHFwgetQieWt8eDLcPYmVCF6AhckwcClD9ZlYYhb1TmIyT4n3I4QoNme+G
byx3mFqBCV6Z/FET0IjfSwQEJjbeiEL2+cPNyUxQuFNpgRESebjKfkoNWm0lP/MA
+m6qNG/f4zw+55r8+RXJ7lGb0jIBPyOqH9o0ah1/7/mqxigYX1OWTN6IJ0XJRfWK
Wv39q1yvgeR1RXvV6swDAyszm1dZ9LPGvZbjSbscQbSj2gr9AoI5kYb11Ju1eNUU
uma094vE19QP802riSHhQJXwTE1obAklgWdnJCdl/z0mnnqOHHzle+2UnrtJIq8y
lfhqNNP04oGaM8PsTLh2ZiHNAxsplH4YHavjMOR2wmtbbgLCt0qSMQFgw6KH3AGH
OxGWoQ69141WyYnNrmzJ92IkqfOO5EcJW2afadmYd2yedvW3z5gTNCI5jurlCmEd
Wf7Bj7UTf/RiQK1cpajwwO/0ldIjacblQ0ePhneJYCgwcTJrVSb05UVokIER6yOI
vTFFuGLsgUYpLlQcu4Qwc4snq0zylXwJiI3F+/ze5hM8suVIjBXNcLxyV388lsRe
WV60PNDz6nriAp2PjFK+O5JUdatCdL0q6Eu2ThlwEfxfkS4NSpGe65O0TqL/Lb2e
QxajTBibYfr4q5qD6yd6rvzycijACT0I1v5CjbseCGTerW2SZzzr7+BLzclHhk+n
vPfPRwo88YwnGld2DjE12MyBE5Dlv1/tOBIwFDyn+Y1Nga7SGw8ohgliSRmcmdR8
NufIlsL+0T02dm6alqDmWqazwb1/7mPhImL+PcwtSWn7/IUd5qcXRXRmY8TkdClN
EwNAi+rqVZSufxFcy5umObkNi400BVmHSOJPYTaD8SqvCn4hUYam9USO4mUbhPgV
tEb1r5To7uK0U1/zonuG3ApAZ84dt1BNA9b3m58A9r0uRhK8gYdMYqogK1/DuzBJ
yIBrE4jrux0FmmTpVxgh41K8wVSxumq5dqXcLZXfxBFHLYfaIdoedSQf9NwRUqy6
TvBuhjfNGwSBg4ul/K+l+c1AXxOopW4k16+4Q0HTrfadOWrteszn3R418ewrPKe1
tKpq9gJy5AUG0dYpXqF1JkMunxse4skPnzMEggUTR/gtNc12f/+snDRykuhlcJ1L
f9yPJGgcQMpHeqzbZBPIe5GW6J+2jL2YE0K1gV8DC0K7dWaT/3MZlXAdj8Uu1I23
kjFmp+QL+FEUOz2fcyGOwnTgP8HB8XuCYIh1MfsuAlkWV814YXKGS6q8ulJoAg6i
77NQPlB7RfbM7t/p98Xh0c3W1YViuWercWAdP3f4zE3aUW64X/FpPPUesqdZ7bqj
TL9cebCr95C+USwpn0b/j+PGJWnuuEauVUIea2UoKL7Ugz6HYNam5uad6k34mmBn
ZLGMN/UMtn3yAboqeoSgdG1U0YT2YO7X3q5Vt64Z49j76xYGqsBhBxMFA8C7XlnZ
XNvQUoBXeJRkFRNRgo0n6+hP2KZ+uaxVM69q+unl9fimuk91bOblRUhJ5hXmJW25
GBEW7v1aixZPwW2g/ngmZAOPgMgUYrszH/xIyM0fux+3Hm5BnFSzmmhjNV7BM5lM
qLaEYnlh3uSM8A2eBDN83E8Dym8RnjAb6rRSRT1bdwtWZyYktPcNeRwKVpaeMgDq
r9ZB/l2ax9GKxqsEAp5rFtXyAdLaoE2B3BIKoKZREmV3EopqftbV3a29CKYMgxuF
80G1tiBRyBUXBb25HklAbJ92DT88L5SqPdlLrYj5LKw2yBJBERSqbg9xGB+P/Djk
VyvswIe13FtuASOao6eptdiO9rjboW9VfLy/xTeejxEWOaduy1LVjjhFpftKhTBP
ytSHkDp70YaMSnmVpK/pOaeBr0nm0pZ9ELII3Ta3FclVVlrbzrX6M3uJyQ77vgeG
bjKSMWGTWyLgw/DTlYZHEnOjIJfHeApwzysqwaIPjYNTNZpBXSO7p4OPD8t2IA0c
CfHTgI7mJsrbsz8L/f0yWVSsjLguumgLqFxsbdhu7cyAno2B6S0xkhVp+PWDmBj6
GXk+iOK+BKTCsNxoP6LbiZ45DrlKS6NcLu55Q/FNdm4Azy/abP/X3FJTJLLV350a
UgvMwA4R8F2ybUHKAONPzztp2hH5Ot3Yip9t0Pa2k1KH5c0S35CQHydQXRK35WdK
p4FVFEArzns/0jvgnaWvfApUx6lpHmEwBw7yP+Qo1RaTVev2YAwK6bJ/UO3ZMi8G
j5tjaM7uNMfiQxVFTFBPL6EyohsFFluEGQObHq0ySJ+5ZwkMGpyZeAab1V0YWWZD
ojLWsm8Rl0StOLp+B/RHRaTnz2SgTB+VQHYJNrmBxYk97DMTah/fDSQjo1iYbfx5
PTJxf/PXsrPTEjJphmO8sC6qs+le99GvxxhI0YAZH4xUElJgJ00W26B48BpwSNgU
F+r6EQWgRBdIKG4UdPo+dPO96oJpwmrlv0q44TZlppOxvNFcELpU0ifxuEzkC8DU
KSaQ+dO78zfmOfOXUW9vW96oj9wS3IHcyDtkXsPZlrtstSE1ytvoAlMoZMdB8B/G
1pQbyILLCE4UeWGd5nU2B3SqFs6Wrtehok9Rs3ryECZ6F6eEhPvKriSwD7mLYuMw
ejHlcFEfEsjLzR4x/GrLLfBr//JWQ93c3x+IdH4HabqbqFtR//oFKAfO2JwUwrjr
htePJOQGs3gZh1kONi6mkh9Qom5svFXgPp0E/4m4CgTwWWwIzLtnPKo1TS77oa3n
u3l84kb4VVhEhyBMFpsFCIVc4CkF5YGrfqdTXTaiq8YERHMaZbkTTEVvW1opC1ML
zsX4T3MzrWPRJMxB0o2xbXHkQLrzPq0sDDe6ihA1ZqPyDdNc6AgVm7i3/e+vnsK+
yg5TJUANZ5St7GySnb06vYzZil6eGqv5SXM3cE4CJ/4G5K9BA2lixpSN19iBJHJi
8Zh/DtWwZ2FUzPJwkRponAmMdhxuQeGPMQessWtU1kytj1tPqz1bhZdu6YX5M02H
LNcL5o6IAXC+ihT0crPe8+gAB+77KuyC58KCBMPzwtKiCKrFrmthmnz5yzh3djfd
vwOSYt/GeNcHT/Zzx8ScskdFvszRIUdV2aQYaZ04oxSA2im4sLEeqrZlcZeVBELP
5gHPD/5L1QSa5ijQyofz4f8UFekHa9mspTqSh31w2B8dXGjg8R/cLbCBko7ikYCr
NlFeQrf1I2+pbXUTepFQr6qbsZdRZYditlQrNI6yidMgESIJxWb1tKjudmGw5ONM
Akbo6E1jELoSZ/zzNHpNDF+HJvqQe+70vBbC0yg1hgMNR+QPBusdXbuYkpUH4S0/
C3bKLNJJh+0eXY+GFPoD5L8RW6Iqk31Od6YEC7piekSbhrKcEOLw46eN/fDaSa8k
c4fmiObsNsFTpsT+sPZy1bSRaQgo4Q99hcTJfC1Q4yulEK3ujPS+lE445Nur/OHU
kkB42oQjHoTI+w1daVOoh0zirwngC9xKg+fNlFtznpNphEwDbg03NWxQc2Os9eh2
j3Tjrdt2it+T9HtT00xNEpjnWdxTg+p63JI75DuVqD2laIkKMg6mZlquszN3G0Gd
AIe9cYTZKtpLSZIP+iwEakeLqzhio+oNwTQOvNXwlevrke+uxOudNGkaxW7XJXBt
5N3sbVJ/hxOAvon0rseDZkEkzTTYnk4/Ar/j0OjE81hByl6nBXKdpn0nxSIn+8z6
1b8e2YftoMg61Yd5pxK5zfYe5oepZ+Ex7OUh7lJfPWBv7FzO6z2t2J3vBCgaBdO8
rtuksJvHTCtuU3vpE5hob3aztFFyeWzTTrgcGUMmw2RQ0BNZxbpE3zS4fNAnA76b
KgIfbqed4lbcaAFyvWQJKuRis57FoGzMWEfAUZoD/fSzJaHUE7dYhvbZsoiY8rjS
XbJSCNYIag12nt+mOR0JT3SGSQMcblF0YRol7JIRcxo4Ep8ldeLhB/goeyUguuUS
GAyLWpHzXJniKryd1tiFj8OHSOH4Kb6qiXAgnXnGiD9QUKH8hs8bk7gMLBvFrqnu
pXlTtje8/pP6QaifBRanaZsSi8T7+QWAsA0lNr1afdCH62n/wQgDrjdWFeSIHhqj
h3HM1PLnWqh/eKKxqReO455MimTgmBr8FpTC74l2n36H5EPDutRl+KAXspPgwNYH
Sbzq9f7aFhnZ0jczW9ffs+jSV/bhMCsL6cqfqwvzwq+u6kXTeeJpya9AAO85oMXu
5h+4uoOOf2NiFpR/YTf6TRf+8rMchfqcbtNWRq9JmOCBIVS5nV1Sv+rCbzpygJUb
c4b5a2jC0gvMO5YcTtxNvR74MkknmhVBc3A+jI1wxbee/qd0Zc2RX+XfnuhxfeeY
icgqcbkwjDKGplOhml3E9uhLcKOfBkYs29mhavur8uQmI/MQ09W0Sfjrl9M9J4V6
sw2//VWe0z+bCXyUD5t15RtkJKN3+WbPM0vnq3tDRDls1rdDdvlpTWYjPA+ionz+
nFVFoPu+Kb60UM7NOwUEDP3JbEeh3gcId0Q8+G/h941v3H2cj/BSHz9QumbfBF+H
lWc6t/AFJtqlst/8ORv0r7m6kbXYCE0MbvQ32QSKqpkaT3KfYZx27TEWrdb+CjWS
tQ584/GeaZhrfHPFHnUapcdsvFaPnvLL4/WrbdboY62iHqia0XvdDV1TYEgdZTTg
yceOhVnjsl+0zk2PUxN8a8SLZ1myWminUjsS40Jsp8DkTNrX52XxkjSIzVkKlgIB
pN1QI2S/khbRgibwArnor8goBGneggiGUROxhNILJ1IsvNdKABkUgaTDl6mLwyMJ
fuH+dCZm0NW3XS4GmsSLhp3vSRSy8Uuyw5x2r6DKPXsK5qcBpflWJD8/c1Jxn/fI
C/4hjrFF/cra9yxCCJjjjVJ/2hbLgh7EX7jsqEtr01CIJWIWiGn/lPMRw8/wqm+2
cNyi0kF6av76O/FV99zYlJm60Ichr6YPsMR3xVYcF+BjRr4SIcjiyvqMQdglirDP
t7aWFS4HuUaYWGwPoD5cXvrQBg82FpvUuK3FRYA+myq4We967Z2J+MkLO+7SifHc
eqsSmi9M68GI2dRfoqYfEJDR/niUYnIy774cd/8/encVc7HJqMiwuDj62C1Fmz/1
hX+81z5b9Ahhag5o/skH9/gW5fhQd8xQgcUdwMtrtm9D9m15Dem8EXOIpTCGPyQh
eOg2o8U/LsA+sv8Crlo5x1+b/lvEhMeZzlN2G+b+kaIrbjWIYwsiPmwYSqk26MpJ
SoGFsGC6NnffUPX27jXXZUvRq5iQUFUxb2PfOv33NBP4BhkL7SEf052L6OZhU9jf
MWNQB/MsAeyooh4L/fVfZYE6G7ttkpckiEhxUkcfbQd56j3626ppib6lYY8eUX0f
ZNWKAhOhpPjI7hX4cMiWGjjn6KTeBN2R4wZZYgb2iR3NAW6hIqVfdSeIv/meM/H8
6xjyF6+Bjxs3DRz/d/5vJRQJ8XHT9um7nNYm4e2aQnZIkx1hEdmh9vvfaQiFUKCT
8TzNu+G6IxavGJey5yJL9Wd7GxhuTD/TUAAJeeXUgzKBkCaYHuCec45Mb8u+pKBj
gtU/J5IvzwGaUWWpvAnR5drS3lkXM29cQkQFiTxKVZAQIdRx8TnrFv5ZqwTxT3ab
aJ1z5DHNYeG/veFSBtUSPZhSdTw64skz6GJDzZTXUE/LA5UCtJnoCySsN98/aDNl
ldyfh3eT3UNQ1f2l2myftBmRvp5lhv6+3g8CwNqIM0SxRRfPPMgTU3uhWNQGd2Ip
PBf+S5ZS4kerNkOkaFJLef+Us4FADqnxzpJRi9uBKuOVxhSyb/4kQMDgJfBhh3o5
WBQzoBpkDZaZu8nRu+zVnWkvjtMgVAz9AMZ4xsYIGTa5VYJ+NHf++m1TSu+N5335
FrKzWnAz5zxihizlnYgddU6qVBCLp/Cn5gJohdj15HsJThUzWjcx3H7/6sAxUYYg
Ki2lCyc5xOUESE9KpMm7p+Q/zr/hk3UkCL5Y9Q9bO7fKo0KlHwiyf3w+eSzGca7w
tO7sxA2LxCNNaNouIzm9h8tgmgoDHTlLU9Gr6ge945k6y8xb4MvjpDUUaT7CX2n6
TVxkzlDuZbIVaiDYToq0re17oF+gdFxO8cdTBXbujVz8TI+MZ2edI/el64VkVwcM
M4+Xrt2XU+DgJAlueh9aldUSFmmc/EQSsw96tANyn8fX8ngYThZcdjLEQ1vrohtV
fXkLmR+t4LbTM8K/q8LvOrNFG+4e+7ugGOgBzqpY7nRQyPg7MwiI4L7SRGjgbjvK
5+qT9k9+TvKfuRD+TYSJVVtoqLZmDPDefbV4n7BVt8K75yYECzCnOkEIanMSwY9Y
B+fHCCNkW+/d5rkCHgBMJOLwmJTbzOi+nDO9RGiR5f3TyGp46TySnxwfln+ZaTLG
bpaavBYGKTch19kG7/+Gis6EmNZMM2PeWDHxof2Q3QCIQHf60EXbDgOzsjOloZBq
nNl3JdWd5X7JkUTVzIO25EYQRhag7xCf+8osiwXB141eXHrBXn0E1gcoX0VLa9Ro
R00mUeeryQ+TRSOn2Emi213YNmpqJIlzh1OqwpUf+5YJ+r8mekZ8dvhDyMHxZoJ/
KiSoN9+5WE4NbflFF/eyRyvhOB7rng4MjFlcOSS98x9OWdzntktfcUX8G8u6/1us
/pLB0ZCMt/6CNKdcpUr+01DqzG/4VX+gnwexp7i5n+SLalQO28RaefoAG284808A
XYIkiw5rECMjHg9+tx1bnqjGqZI06MPV2uWfkv8VOsjyoH7RH1U+chjApA06xx9e
SwDDmnPuc+0ucybbXd16nW0UhHOAzVv5jfgvOMFBuUMgu8AwsDvxAPOsMge4BkD2
LdiOUuUHyTGdyaF12WBVCireIXxaAZ6dLd6xr50ir857ODrXQjCANe/sTnjlEafu
K1JxOZkv89xWEAVYiY2UTNhznJwlXvjmzE6Eb1lv/ogvMBay+9NISJF1pXyJa+rH
kdlilOTk1g4vZa6St9ZEy/BwMJ1/HXNpGTY7uoGzEa77X2duw/ALhqZr4TEpC5ik
hBZp5nEYQG3iH9obwKbIK1BDF0VSI2POxxvflvR+mVMILXIT7/J44mbtGHTCj5Y8
12R+7Vp5uPS+VgO0dnATrWXSB2tzF66p/gsEr7m5YlK2Y89slYchfoEuYarQAP2K
Ccm4PJw+H8JL2uKYtj+JkTNTji4JqPZrTakZax2YPRYpRAw9mKNfWFlAMRmCHBAQ
4xc5MTLxPZEi89xr/YOrzLQxwkLyRi/EXcsVcu6FQB+Kg0CSCcQ0l9B+4qBQvNF1
5wsV5QNAVSnLj1m81qt5gxLRYaPihwSw3WVsgFW4ucOqaz6Vn1fHpyEtCVT4ggMi
4RlxGjBYUp1uT9unbE4/UCoWqOoVI32l9+AP6BRwJKMhPszCik4sJdbcJkOayEHk
4hEF92Kcx3oKqwCy2px/JDILjt9i7WH/JuPB1yrddTVrCaywt3DHZvwcWvQTKks2
L9HBldjxC5oUND1AJ4jT6yFk7kitGon+HqkUbxTTTOSrlvTkB3uHJu68Go0WZYKq
VVknmYy1ystjDQbngU8uOkQQKXWCqUhlwk66ZmwRC7fb6JC1powz2rKesLabJfjc
ADuQah46vj1kgO7nubXGFifEGv2uuvM6XrJbi8Tzy/RrBUEVIKJbjY7bzJ2kIxT+
C+D5sZWos1b3FqnEmGg8CFLkiR6WzjLsCVyqtWREZJC2b10U9rjELVqkT9AcpCtJ
op2x/jDWh0Sj7KUYoXl63QTF/5Do4uJ34mm+PzmGMCS6LpSpqcvMb8wp5RIaRgfN
sdZDIRXB1nbwnx0zrFbIUTUgiceRW4FvViNmPqheoEZbDb78s32k62pUTc5uuavj
iF7TBxyFkgU5OSAtXldiq94ITLY3Fbo5/n8zqU33NlbNPHpLFFeegafAa0juPau5
bRwPHS7bFd76AaOGRkQdyEddVLkD0AXYneFnGKfrL+9CRqYRfkRs9Cby/3yMq2Ov
sa/6ivEzvsO/b39Ql5gmsXB4XGEjc2w71u7/ubOTiciYUfaAco4NKd2wU7ccn1cJ
piGRWE2ZINsPzgC1SWGQUlsjvsl/bAh353SW0RTEBescOAQurym124Y4YBFbFc+r
mGLjvM+9UEP2DHfGVJ7pEdwKVjXDIU9fTrBUpJfW08neloizTwSAB8JOeztu91GQ
m3zJrITAE4KubiSJEwDzxsjPq7NEXKNJgBXFbXj+FYWr2SYtcyrvk6vXf2tFh60+
STuVwIlKM+98TUWNsmr8H7ozwbfY3D2gxuRe1CJ5LI26vAHUdTwMhfvd9A4JxIII
mLdPZsmpwFAoFoSkdU1hQI8fwEuzD3iDEp+x3g3StZPr1KrSZAzhFfYRmDOtA45S
6y3pZX3KA7kMPkMaaT/HpletbH2SjTedj7jrO3wgvD2MU281qfImGBDo/LphSkiP
vJu3/mZ0yueWlQJoR55v4f7i+sMh6Q4wkBoKrFiVBssk6pNL/xF2WwKq2FoeszR5
gcgm4UrSis/m2u5xUpRWFt++2ZLlMLkj3bdO9ZzyMdUUBpfyNZh0I1xbyUzMKigZ
evbyYPY6cP+mmzw3jKzrtkKR0DZWoNHfm3lodswfFgsCgpIvrHsQgwrokDtRz7nH
IWtMy1MO53fF4AzdebZmjZKbdm0iJYcpel/k2E194RLZRAYk+T1q1Ll73022tFYc
gEfftbAx7uFYGYIadjcuA49tpmxM2dd2wsSHAsB8gPt/2tD/f4EH0pvquaARn5S0
TPoCcLSJlYbW7w/+n3DTBT06RbVZNSrCayZWSawJhTuAwNMd+FmgE2CmqFYZM3sH
grbZOfRhk/J2uytlgkyg/763p/RkOGfOZ+R6R03+rFOTu/9wSiG7FsHI0N5Wzjbk
BK4Gaw3tZwLQji2r1/p2VPlyQC93nzCNfCxijmfhrAR7U/McONrLG2/IFmJPIQI1
CZFasJH8HpziwD5ktGgyEN+sOM5laoZCB2bGsZwiBssXE2iYQTU9hF9W/Zpc0oCJ
VyuMJFZXOEoKPBjJeqzVz9bn+AmoPPq1f7j7MTv7ElNzx2xCslPs2IFe5ow8KYfz
fFWX5h1CEpFy/f5L6P1CsCNcXcNx1i7p/UFuTACX2xoG4r4NZkW+adH51QxACs3V
sADPuDQhnQP2g/AbinTNBdmxpq9FNzJWNkJMd4KB84yOPIzFW55oOc1bXzMnSnAR
L7T0V7q0iuyz/cwLXOnN4FbCHOfacMjk1hOV+5pbUKlGo2ravur6G4YmnDaDSkZR
SiV2GBqnVtY2Uqd+4A8rE19LM1WNx+cLV+qJMnyqSkG9wzco9oE9LrVRYrGiL4D+
u50sO0Ff6yhq20PNjTEkZIZD+rRTLTStVqQ2nV/XW3YNEDsXSXnTDvNHez+Q+cJe
rOoV/zXLd9FHkuMug8q8TeQpbhDUkK8H1m7nBTCBGMI+Cu5Nmtlt4s8x0I8HquPD
REh4FUBM2yGf9t2X0sRwX+74wXQR4JyaTLU1+vNyo0wcgs4yUQYoPehlaLxDJ9Kv
FHCiQDdXcBC9y09szWNhG1qHz2EgSqxqgb5iOWtXTyZLn0SHI+rBs9g/s5mHesKn
HZaWd9SEd8BefV6SwHqFm0e6kjspvZ84vrJHjNVB/pE279ZoJ+3sMM295pJOAzyE
ABSBvZBNck6x+52B7NqjYJtSscyfQmEYTZrY3crsjJ9MHZNo7G6Td0iKRVJUAM6r
saYsra9kwj8QCELaswtjAS46S7GGdwjiVlmVvKdhxdJsQqolJM1JPS2gTwef2vXI
5tElWp619ValiZ5XdbGZERq0OtGVLIo+554sucQ/LesRrf6MibGKNsESXcjS3Cis
gph1ZBKIZVNJjwpkPvYhQBJHP5cDMcq0feo9uRWcfE0ekf9/6jfeBg8rMmAP2UWW
rSSqMWEPFQ04GlgFsk1FaiZiWk4WONIBB+AFvv+i8VG4WgMVJtb/FCg7CVuVmhYr
1TfMa6/fCDk87/lw8mMccTXcdPZ3yRDtX0aYDRjmQVNc0Ng8UMVzWlM+s4UMZ6xa
eoT5bnEsSpn1uQWqvczShmb7zZk/EJt1VcXZ1ASsywhd914ODW9AwRywErZJJaA3
tElI/LBGIv0GVab+9OBZcU6Ipcyoia0mUNxsgbmU2zmgz9a3luHhHzCkzIZbfuvC
njEGkPH90afTC+UhWQyKWdEdlvKOYUaBUpthAy4neAuNJU0sWsiw/71WLBJozmWg
LhJxZeQShVNfwcOmmHvRfBf7lFPomjuLJobKXKaUNnGpmcfuTA2u1eHy0pnAvqsV
LtBou0Vf/9intuHpO1oSHTw7KAsv3rpAW3U8Y8NjVSnWPzyzC12nhs/TRfr6/TRC
dat+gIc7NXW3NcNetqXyZ9qkzve4buPWdD0If8ad2aL7NnACUXwrluUCngY2t7QO
vIR2lrLNl/Sm68QyOcwUYM9JZtWDyGiLSyceUO4fmU/17uDsk4Et7I7Yj0J4/ho4
e3i/lADdObTFFqkIRLgSomTEY0DC6YgLH2YYWXhdlRulJdmEwC2n9yWlCRywYswm
M2FnGWv92tTUL2K6cY0yN8fA0mvgwlRn8LzgA/JGrshN6q6hXi2BQL0mdgD5f0nQ
DsiNLH8HK86sw3E+hL7PrFQmVMqAYmKgPWIoBMPe+juAH0wzHvLxPEd6S0l4euOV
AyQ+K2MEJlhZRc82gg3G4DPZwUeyS8MyfSzBbOrsFcNVkXhyfabxc5t/oEuxlbxy
dsGrS2zqWmkMQn2z82nH3iff4O/H7esncNDwc+i43/Ly5Hj9oKYb0jIPolWtVbfr
sFaP13+HJB/PAUKI9m2SGEG0eBLmZj+lYitUlGt/kYBp4jNR5H8m/7aO5LtemYdo
qhUa8xvcl2vdKCkv56F7jlEGPaPaUNsv9e8I3r40ToaUuC/MoI39cLqwozGoDoX/
ll1moMVZ00+AnyxysUaf9V556iTEYAclU3PXLtNF545iKXTnLrIZpIc6LTOFbynn
ucaNSp8B4gBWKWBRBZHfIp8yAtJqAIKzRYSbZysvQbEnKLP+eL+mOePpj5fIrp9h
D4M59hREWeN6f3/G3qADBwjWiFNjV6+td3qflTTS9DA1rU9Ush9gXK7DkIw2aw1a
VWpKLbNXyRxNPJtRtn9Ldmjy2vMQYp6UhrHJ444BQ6gGE1UJpoj4s+IcSpqBIGrO
v41gz8l7TrfCnIwE+Raffgv36Zu7wgGDfsozMwkyUazJVyUwcf5aguit3SUHPY7Y
cNxmPtISafkR6kgUiPyp0Xd3O2jzAdIDuQTCKoMebeSECSLwvrnPgKsmKR+SZIeu
qNO4yIpuwyHOoBemf+MuRa/hzEEWSQ8QB0l5fML9Os7R0I6vrp49xYXLZ+yWw9RX
Zgy1NGFglC2IZaHc2ZMh7CqQjQikB98+mnMBSVpOW47Ue/ltVw1cNF5PYGeuqL1x
OAfoNFmjelgYk+oMvbEkVUvclOtcUW8HScyKfs/tDI4LZnXIvz9EGq5Yuw/mPQG4
9HECQ1vUqnPlYO16JtuhBlQMm3StdLGMsfpDwZNU7GsnG9skbAYqkbbYhZohv0nL
SDJCUC2dy63PoohkHVZZ8WbbZt7DclBjB8mX1kteEJmeoeS/EM7U0qDbCM18GUah
XQgYxoDM4E7hyrxZUBOj5gRKvnDVQsrH8X/FdFLeKwZpJr3eCEjRBmoPEGKIF29G
IBYRr4mYp6JEIZ4Zj3Ml4IOcsIfmG03u7Fu93O7jnz8G5BXANtpxN6XFFo/V1PT0
PQyn7pdvDY6xHslolfi3vV3N82jDJLzwQj0AEeZokDY4QCUGSR9lmxVBttPESZFq
76sGfVK2AJcSFqhsRa6k/LO5PJzZHuKSA4VPFStJ0Gg4WdhfLDgnolzIfjhm6tqU
/Em5xcgzMDMaI9GKNmHc+EE8CU3D8g687ZeGrMUDr+Ewrhm4yrcPvhrVA5cVOPOc
bLqr6DKjWg0He0sWVg3TXdRdHrc6rg7gg1felNkMzXFlvpirR67mhm0pHu0yXUqq
dy3VwdobneAV+AFfZDy8LadATQeJqYpNbc5XApb4ynlO63zuJVJ250xAr3rM5peb
ifwv+yNNDhghlXexlBtLQg4WgIN5fekLTZ2Iv0EKKb62dtBKWMBYXrx3qikgNNdv
MEvA+yXQMjpY4PnD+NCKIo0MC9kpX8y9/PNw0bYn7t1RYMfbk8TiLWEfOcXg8naz
cZbYR3QxeMTTTtLzFJ2EOISNJ1gkkCYbBPuA6X+pSnyjGJJvv4zVm/GjbeW6C904
oLCn6BQ2oGYpqJlS0MO8pBa6NiIxMr6Y3MdVW+QvkcT/WHSmqSo4+qlVNh7QJ3T5
gETYd+4a017Jj+rMgu9ZGT26WiRpnEmwbUJaoPNJzZ5QDiFBKirG++MzvVovreP0
jYkmaNTdcGWYGMQ+kLUYyD+C1MYXNQ15DKQ9qKyMkkzo2usFdG8TfitiKx1+BI/x
LD9t03St+1BO8HGGPs7SAAb+4XBbHBzaXF7F6JxBG+RCO8wqLXnqRfalKw9XhCed
qUs9bY5o9xLp8mWksrzYa7xxRS3rgjBdYL6YfCMonjayWZ4Y30TSZ0q5jYpXgUAN
4jyUs74bG03qPzXUR+6uoGRSuzOsYTL4lH5BxJNqGHBjxteM3PTyMPgu/bV8N16T
JH6YAgQSXCa/EMB3wuQ0WungsUJFKQ+hxk5Fxlxo18DUwgaPZXsX1zf0gSuuKpW+
12xYUIwUj80nHahxqmAnGtNltUsuwaoKWiWefB92+l50rikSkApY69noBbCmajeM
TD7pgntH20U23mbXRwsqZQ51UuR216Hc7lBnBo7Ed3EQ7B5ApLYhlew87PQ7YzS2
TmimF8Mxhprf+/WDP0TxL8Gj3dIkfILQsG2SnZGa0JCIDoeDw/N2lKgPFDoUMQj+
rgbl2XatXg7JqAz+H9y7Whgp8uZbrRaFCRREUR3zwFYYRmrjDMl4yBCfeSbZhAza
MFa5f0N0PEm/AhTFVPBXgGdLnSBTCY4dPnbY+iEEBsQ00fDl1QymnTyrs+9Rd1b7
thI/F+kwmU8Hdhl5ET9YyJmL+WvI/jBa+ng6ByfxjxuqGW52LipVItqZhzVNeXLS
LRs8JYOD7tB7dsFYBt3k2njyXV5CiKul0lLSg523GfJU+0B2n9ONOE71rvNaMtHb
O3NCWaGtP48Oo2JkeZEeUJYL9p03lQQqhpOy7kPKhQGhSLwMl8np2UaVL3B1AyuQ
yHwtiD3QOmzXv0VZ6uKKuTuCiTlUwMz5YWcM7wCznsPLHLdI7mC9uF1aCWz+RpAE
INTHvm3E1c8yRfDzIhBwirUPQZtBsYxlKVSekJFo9N3pD3kfTy0VNjrq2jAVTJDR
ArPY3d6pmUwphJauki9DK+8Ak73rLRJuEwVopGfsa7izwFkhiGDKsPJ4p7XE+VK4
bFjPmnkMrr/HBDBUfbpK5aXiCOtHJ7LYe5dt+fJwARpz47l91uWLU3kAd7UQA2xc
xKpOmb6WgezFbI97ghqrTdOzBldcmAVLJoGUsqjhwsluc5Fkx7QotE1NeVYVGGok
aCh+zujgd4meaKZL0HWQNcI55eTdGJMFlE9BUNIlrNxWxQLiA+TPmhfIYjBwfZWd
1V7If1hu1QyJgUXDeCZQWsPfRdlNJPOyz5eSY4w/chj2Wcmlu3f1kTlVNIbL5dHU
+tAI/0f9C8yKDBba1kAX/7FLF/HqJfnw78LNMi+FNRWrvlHxWVcOQM0JvCo6Sqp4
7FcofFhEP2b8IhXVM4SQ/n/8Mp05h7v+IhFj8SFFU74ICrJvCmCi3LY7pPMzTOfS
ljrAp7fAm8nX0MPoAkKb6AIcQOOtNaLP2wlZW2lONig9BdmsF7Sfo6lSbVrkWsQZ
Rk2b1EjwyF0El3eTzVPjSMwwX9FKSW9HMCb69bb95tYDciB63NGkC4aPadOy531K
/H3X+QnzHfJOFYrHOVjWwEEcL4W3R/G6qR7iLsiMaVZ4tb16hENXwErMTIwkP4PW
Dkg0tDDPzgK6kR/dfFVzG6vDPU36RCM/SxscqtJkM2dLMhsqqdfuF9hNc2zzvBut
Bd64eEhX46srtVk31McgfoP/Dtjw1sLpJhhOjb3flEM1jzRcvX0tFzYrqfYYAyVk
0m34ySqBcDDtj3OAm/XQNqwnQ/D+1fub5W29oSm/+pE2Vhs04sfbnw0egReeNfhv
QrOX3E1DWYv6/JuGTpIncX/AWsQDktdNdQfk83TckRoxnhxosZOfL38Bw6K3sK00
e0CLnewvAsGdR4IN7V3p3gjlIAX7gnIgUTG7vir5VEPKfBz/fM7CzfL0rTxmUyfz
qPYULRwkQYHH1AJSNuU73/qrsDDl9G0TrItEs74Bfm0Ebb/Xy7qrW6Eawgji+axH
0sIwlgIdg2KpH7wxggZDWXJojBQCHpL3zDMUn/F5/0x3vfLRvhYZijkphxABDPdZ
RkeXFxR09F6xw5yd/r51JGTa9Omh4UOZ9C7HOqQAYMbMjN4ex1vzKWF2beVTqglW
THmT3n2ZAaWpG2uKSEaN3B9zRKNTT7bLcZqLTOWuo4agAI/SIoPqrX4yCPO4L6Wc
OiKALyKhPiyqvdEGrVS+YAc/dgm3tQEG0Hbu0N8ukSGLvGA0vQwoTCZJazjGMD6j
H2vXwWuvyvFv+l+N54svlmVhq0WwlmEjg6hpdDL69+x4e+QLL1+PQpcSA5oSphIP
12Cgz6s9mn7J93iAlh3jQCKVqhbFsE4P16HzMYlANwDbIszD22ewLmDZ7XukfIlw
67BnpcioApmgp8KskIb0apf2yA1b2vo2MZtjFLMI+P0S6lNXCU0tiVzUpVuUGyUB
+SQMfeYb4sRsQu+prVj/3QLutzCPP95tXn1sx/bjDAvzVAVGWgisiHFExVZtdMBT
SVfvQWGzM2itGIa9o+3s589jwMkRTDBIfcvDfRWqLxc5/7D4gfCfuZIRQHg/bDvy
dpHCet62lqNeeV9zJ7ivI+hadb6wo6wrAyt7WVKiNggP+WinRYUfQoyGJCL4gZ8v
oskrKJqtYezBfcrwBBqBVZ6m6TudG25QZkLv6MrIemrvh663XKQApuZkq+44EpDh
vld5pl+5LvRWm9L7WS9uQHEAYt68X0GoPxytIfp25LEnkCq0xqECx0fe3ywZnALT
EUZF9ygpVSEg3tCVcUAHOuCOsnbKlk/qWnKrWUjAyJBq093rZGSJ1oMKWMcSGNwC
4ocW0njNUNlx/S8f9wyt/vqykjMo826+Gn20mEsIsSZ9PPycBJI6FBl/ekAItd11
/Lj0ELYFAWjX5Qun90UM5LYK9ny7gUsaNeeGLdFJp2oX6oxhEWT5mXlc1O4qbWNf
AhtSW/LysfAI/tusum/CBEl/W8V1tR20gVjcfv9SSVX4Fbi6lSBGT1l7FX17BZ8I
vFzMJmHxCtE/HtXA741HlDl+xjiJXYjavzOBHcuY5IPAgSVnuQjyt99eprh7B5Xu
HBsI1r9Yyfm98MskVM6YDCRdT2x1CT59X8laK9VPPCjDx9jgZ4w2at3sfClf/5IV
OPz4CVsZvtVNDEBMf3SKVLr9s1OPQpn66KGOFokpfrzIAakWwhGFmOJ/nfxaCcI+
83bAY6xg/2AX8XMglAPkG/zCk7mSO0gxV0bDDOA5c2wl7vY3DBd7aH04IojJy7z9
fOpyK2O1HRTsBJ85oXFaigsEZ0XILo+iw4t0bPuY/4euwu9x7KUbc1FtSgSO7/GA
N3gOjZXAsuESVmh8LpDvZIwyT0/xvB+8GgkrD+XJoWC9Q0BznXe7J+QxShsIBqgE
A7w82gF0Io4d4rKkBD7m5Kxh9N3ndiEqDSoPYFi0SYQuRIUb0RLcwnxwuA6GfTAJ
/6p4QLaToAcl1PI32Au48FftvDK83GhyJSSrmxUJyWAKzvylsuFKZmqmZN3o6xoq
e+O7OmXdfAVzQb47npCrxLdKd3jMZsHEKIez9kibIqhxb0IbWEg0J7eh+cwuSEh5
I/qBi5PpkU7l0I6s5u51+9KxVJW/W6CuaTb8C8ZrBiRFRsD5DclVI3/KVq3/wNhv
+0KY9HcQdRXzDwY/F96pejWPdSv/44JOvSbyQTVietjKQ2dfTT9MoTeXqFjePzFK
e0UED1nuR1IWQ2Qu4v0yOUotmtULucO7Dc2zgm5Goz1d4HdnVfA+vNpTzMVL3Zi7
0vDh3S1L1jS4wgYvAffqjnDlyer1enWBMD4dU1IthlngMSp46yFCNf9M9Zqpe+ZE
GjAOxRl+nGbqzCcr379kxOGLMLz8bZD7d73q3sh9fKZ7ynhL88JEea9ymE8Ta9Ah
mopGQP5U08xbqkbKUuESt9eFtYCIew3lKDsluwvG5/hNLYF4vymlR+XB4tQKpZMR
NnY2oTATkeJp6h4gPXN5Wgz76x9MsS3R1T3FqPRQflpq6qxK8BbwPxQHT0j3VE6K
2EfXeUml+7NtHhIogdhyr0g4YVLHeS31UwZoOZYQlkLg8L6YyQzICPFReRR7S6mx
RQN9m7gmiq3E953w6JLm3dI6nLjR6ve4uKZ8XkBSHQth0y4hGiKu2uTPnvLBokqI
FQgl7IQdZCQ85roxtHmWnwueOEYY5W8SuechfuNxY83j2UwF9P/IpOtw2LN3eHb9
lS17HZojNmlHT87dkFxPrM3lDvig0kSVMIJqsfQjH/EsdmiMrsp+sCOlfPyS9CLo
MaPvAXm79sijU41uKLYs0YETCZGsDJwuqv9xhNDl4onlMB+zCCrWBroCXAt7daRj
I0oCllwGrXhcn3N8BFpQQkgRlt05P9nkcDfaAUPHalFQ59p2spOy5IyoadDJtKgM
61JytPvJCxGrqmNAtOC2/8O+NiURbcvInz3Js4yu8XX8TPIEhnYh6myMXMApZdQP
HTh/n2I3fG43myGyHtpIWid0saGTLS2uAby3kAfvlYWJqha5y1WPZA3V9/tyfzvk
oabDkl09LHZEiodeU+qLv4UO9gx3Pa3bQ8h7Rx6u+D8Yk39atK/To2XdRi49Pkfw
rGrIY55nRg0mXxAoxaNu5wQmOYZ+WqpZ3iHV7TH98z8GIOpZZ/g1zKoH4Obb60CS
n8lq2/rbdet2VYXVCaanwXpJt3kw7kj3JEsWoVLOe0rTjDjIp4GAmj9E12Amr0Fe
L104i4jnP/LUxdhdTnY429sapr01URYyt5Wv7ELwY2K/1cTXV9Z03Vmhs9UA7AJI
wH+WR+2EiPGuQw/6v/b+1TAQ8KX8Y9k4bQDN7ReWvBGFFRNdRci6MGWaB3v1iGAK
jrzbJ1d7GHNmYrWQBnWNIALvUcdP0Gkulsgz81p/odurCtcPMVrz6vpOXWLdpGE4
dMTuTMhL0bL0+NlsCq7ZXTLyKfZsIfO+ebO/cF1lKLazSU9YU+t4jM+ANXjY88Ao
gSLkPhHesIzR6r7bvG4wxrcJO5QDeis2dezFQ9KuSE76B7nKSw6GzmIhYFf2JhsK
YuyMtaDEXLCjfURurkKgIzEr6oMoFVMvTUa6rLrbFOCG1abcIAiHDACbSHptbMm2
+vHold6gZwDRzSujPfp5FIOr8V4DvuABB4PWhTfjRTwo4RjumarjYJ61nqZ1clPZ
TJ5qyJpyXon2HrTUUe9fU3guVS8Pz3fVP9fM07cK9zwNPl6JqrhjHjJvXcQMXTbU
/oztKdepSMVj94T/Hu62G/vWIRqXhWteuwXRUoqy16ygjK7kiC70AXO+/0n3yc2G
kmoCQObvpjU+H61ndvnVSzr9bbLxq2emQiG31+t5xEf5ARJ+laHwKTN4fjE4IDWq
SMp9htAvbKGYSEpNT8Xths2rDVmPVeBGX+OPA8EpvPQZwdhc4RWf0PAv4v9EKv4p
8VaKvpB36vWJ/l3PRKNtQURdO9OuGU4gx0wdgTZqcSdkKaEmO3N17KTkMHi12LBu
Qj20tz6HM3GGZpzzzbWLQ1K8j8I4fg6hPrV8y9LczOP9nUZeEX3Wb4VgV5Fb7JmY
weAq+LlRfdZKdSsDqZI/lj5DzNfL/bhLbXNiNSMmqGWJ+JBDyJAOytSVX1t8LNaB
CsfTMi6i5v+HByZEwU81fzWhzsGmYzKsSGWdRcl6msIHew3UrTUXwGEQfQTtjZyM
QvfAEasqrOTGl3N+nS07bhB/IoBmjMLAL3iDoMgr19OrPtmMvxiu4wRHdUDu3gqp
wU+dLh6jSknFkcEo+zvWPNbdkd8dk/grrWkdzP2ETgrYkI5IrlI3UQ4IHHKyq8I7
8E+E1lS21Efth7KP485XD1LqIBq4DNZeXtgdTQbPMzuMxsWjVaSJJC2b0WuZDFxG
mHhKZ3iHml4wTf4F+exv59l/i26PbX1b1X2fh23HRjHRbOYGQKZNKSYdNiNDiBeW
O51+3OYPJWY11naBKXbLnaw5b0+4ti+zk8eZ6nBMLAmanmIb0ReC5nYkZE3zpFGV
yvvhOdqq/m4mulF7olB8hZ4Urgrz3jz57gtNA45HsWhJ0idcNmzwCQ1HUm/qFBA9
kdGKxl2XmoW4CEkMTSAG91aQZnyJzs4quWf4p2TQFWlqUfq9OjkxrHjcav7gQdjT
RQmjWyd3YNsMcsPpZfLllTU76IEZikN7dSlTolKnvckyW4Rf0aREi/8kRQXqbBPx
ysMtA3NkaO21Br14CRA1Ia9pCebhMDRjMR4KzPSGJ5+dFVgT8l3m6xsJ8entzj/M
ME6qVvmC1lVGvDP7TPNlBhw4RvJ+HL8z4pLZi+xH3VEMOajkOm6tTBH1/944uAXe
NuOfvleIcLgtsyX4vsQVfVEmmmuVY26Wi7VjLtDNRqzH+TDEdD6ePNKsHiYj+leH
rEl9x2eA00qKjXbjhyc6tPi1WubUevCE7skcUK6qf6Jw0DbHmpU0JSDyBHVCmhvH
hgfkNlv4t3GVhdNxrObHdjOWvV0ATUL88izj1/Eol7s=
`protect END_PROTECTED
