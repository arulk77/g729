`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBox47yWnJjGkiKW0LYhmIxVc0yNjR6CZILPIhGXp/Xe
e7fel8zkSxufLVrPLw1zmIWA6zCW1wScQuY5YdVRMO2xqo4q323g69PvflLfPknI
ZDVMmrI2QljgQCcm91KwOfkiWteLH64SuIC7dU7h2AIr5H/QG2aziNnS1VmnLLoS
9CKIpna8Yhz9Rflppp62ffQ/1TuszSOr8JIds78RqprDRwkj++qugrFP5jqG19p8
bGZwO3RGvwz77rMYhpurGFpnxGG3o7hUh6+ViZfOAZIp75ogVFY3SUFCIvgZbqpX
WOztMa7SOYqkqBbHqELr6SWjH7KGb4RiuDzkrd/VQagsXGpNhwwQmFM+e6P+5JAh
mXmZ9sdrvaGTtkLnvP/S4BV1dlH0FTEZdcwuW97SEuVBnvM7RMuNtWJIHDeciNq3
SOnMTrFvhtiJf/PVgmhOyxEwQWlGp/rYlt+0+pOlij1IYsGA+ihg6CZTtKDwWK/G
`protect END_PROTECTED
