`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKVOrMz5H6YBNVnARm1VLGB+ptljoJvqtwdw6rwT8oZj
PmuK7vZN1C4c48H1ln2VGxFwSrIqqQciXzn7JYEfGLenWr4b9azvyqPnA/7UhrZD
+pAfXujEnV2a99VEdwDSQ86He0DKz511Q+Kwa3jxQ7AtynNf8UYhEiP99rZ82cxv
cUoyrBh3+NzgKqqHEVPQsqAyHwyRSy/gce4aNnKyNsnS4fAKjCddSIZ3I16+Rbsl
PuPRIE1Xl5AbRn2/CVUJP2UANUoYY4wHZ8Mzhn6V2A7GoeFoE0sc8OXZybVFgfvj
ypleikvI+X8uAD7evBosB006kES1taeS9ViWBn4k1CfflZ3khYSETT3iNmPKad5D
MD8VocA0mtXITQsvYulzIqWeMP1GJ87Cd22DlcJmpV2TAECy0tRX6gPgixRQrOHt
5J0Y826N3CMYWeolJx7wy3ZzXjCtXdwecfBoEJz28HqOHxLFvprUnfuu6aoIDbzg
Ve5g3od9mgonKz5hyHKVbQF6ieToKA3EAjTKS2/wpaI3BoXmOv0fSMjM6bmE0yRD
`protect END_PROTECTED
