`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxLMECoJDla1Mf5ZmADwZcth2kHoBT4aV4nzGvBF9Ftd
MARa5Tuib0YG+DV4P7TjxMuk40g5HdkIKiyx9bHsj5yWhPUCcEzxNAfuXchSnehG
KaflRX98QQBLna07GVFQ+4y0K1MXamnBE2AfnIL/XQrih6sm9F+UxwMySflajdX5
YGvtKSJP3aVySfjkgn9KqVW6iJ8EPNFbgKcs0DfMpuWkXN3zsqmPLMH3jso8EEEj
`protect END_PROTECTED
