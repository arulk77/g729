`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKsNue1sGoi24q2pZyFiK9PEdkWz4aqfS4J23uERgcUQ
nnmq123x+2f5+pWzzsEWpGLKbWXIxXjHVGC04lGlVz1d0FvnIt5BDvh0kB7l+Cio
9Ey+ds3nhRtHayznFvMn5boWXe5taeo1vVs26EwK8Hf+ZyhgwCo3heurV07v4J0n
13PhODTkib8zyoBS3gaS8CpWq8RPQRBBQ1QOeIfsDCe7cLc1VPk6WeZo5Cb3B81q
L/2VTAZk+LVpHBZf99VXeLEn+YWumbFJfMjF+ng2/E5n9kuahz0Fc+y08bYELQlE
CHpaHgn9QBgBU0ztQlvydyC85V2Jw7Jv88ivcnPcBqs/K2sW6U0pdZysUOQyKCgA
AMFswcoHGGMzKQcVzuMog3NeNVeq0k4f9BYghENs87Mdpjg4RYLQpRF8aEBvOnkE
48czcWWcJj2hvF4EeoKutaRVRGaCwE4EY+zjPieBGl8=
`protect END_PROTECTED
