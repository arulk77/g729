`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42F5LJrZdE16ZvAJD4xP8MPB8OFyTHERjq9h32kYmZsT
2Ybh5jAJlqmfiDQvOTPUWx3W8haCwsSAP0sspMPODpwKEmOJtdKFs7OtPSN+cCTB
wdoAEKA52gSZTwyKkr0lTjNys6TfwsyyhjWjtsx58FFi6ndcPgqawIXf4JaFl5RL
XNsn2Hd/SRRahhtN6g68cnz2dQvS+t4/DdOJBORBjcYO1JodSXlrI/V5oWy/dPij
pXmIfFRRRx3YEgTa+C+wSiTdWCSU3+JsH7xpJI7IqkM=
`protect END_PROTECTED
