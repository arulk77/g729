`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveASrUagIzA0LVIxYxbJj5ModKevbShNE3qrG5tOkHEcc
jZT5WC0ZeBnPfMqqwa53RfH9ZZmT37/r9s7KNih1nz4MFCX7gXGVImKxdXpo+/w9
vATxwbNfknl+Jq1dCuNpEKmSTzXd4gIkUmecBKOJ1yQAI+R/1Jast5+A+yCObhjQ
DtNrRwwTiNkH+cP11mOoZhrKQMCRqoN+1AD8EEd5312hIMORC9FWNUSr/sJlxfxC
`protect END_PROTECTED
