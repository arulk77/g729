`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLjUSJx36IdlVb+xAClIiH/G+lIx27cBotQaARdQIVvz
VQuYwwnpgSFPvnpQZ+ApsA58dMM5boFiFRlqI67/Iwn6P088NXH2hE3fNh3XuYCF
d0rRYTEYeIFBXWqE0lVM+3JHkN8HZGvqu+tSy8lT0lXE8kI/gvF3vcmesO6AbQ/W
MX6vO07XIJTKcQplNbfgTQ==
`protect END_PROTECTED
