`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xhfiCBtIb08qa6OSgG2OdQBNnhb6wQ+ws8Vs0mBKgmZ
3bRcRBv230hyf/a80fYY5VXiiwGAzqABmYYDTrt2wuDxQPMzOCQHbHtwoTHSpJqa
FCiGiOgZ3DdeaHvARb1yGDnv7UVwfgbXbCXX8/TXbl/gAXlW93VQEuCUExXJUPo1
4NNBK2UdFfwU11Y+fNoXCXVYYJk0ljBFhFo1Y14Zc/sPe193CO86MBEblVi+NaTj
WFYfjvJ4DLEDnfOFAkbvIxMeZHlqDDZD14vt8/P5WL60WSGD8CnBQQkwW99haVSf
+UmQsJzW2rhlBKQmuz2kvA==
`protect END_PROTECTED
