`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/hzqT3wYM6pYgCVJGtHQceZkuLgre+WfB7uzpuLln1dI7kHOyTELH146BZ8nG5vF
3aoI1HQdR/1sj2FLQQoSxxHfF+OXW7EAmxijOsXRrV9VAf8Q+94BCS/ZPg0UTteY
oMcwcNZ3J01RT+lzoHJ847uPHWuQfZJsl8LuqyQXSnypxlbzudI/c6TGeC83T6vd
03Sf3Kf0yU0CET8BogYfme/PdywPCURzZk+97Ps2gVA=
`protect END_PROTECTED
