`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7Ox/Ea38rv35V2SX8rLVt5xhdqJ3V8s5n4ea0cxQQNyB3u7Y7evfwQO3IQgdvoZp
SMtrGst/RaMNZX6JR85UucRWmLe9i9B1fdl286qTINOAop5yBYm3vj3ufD5Mwp0L
t21wkGbfveJGf65qTkXtWTHWFeWeBat9cWq7712ayfOOSmjJzz/ya522YyFrgngk
yBFa+UWSrL8cAVYrB9VCTZ01nPMm5jOoxeltF6WlR/2AUaViUesHMVyoks5au/Nj
awW1ktI1+4OL9I+g3XkwIBnCMhf7NruzhKOKyOg30dNYNPwAtKLW5TjwSAELY0xU
0ce0nGecvugLWbBRC/1KjKgqiEln1aynnP+YT8DWI07Cmdr0INbbicIFbHi+ONR7
T4YqJPtbE0nqyrezs4lnYgjVfKc3MomkVA/HJS0vrLxZ0EAqO4pmlqzjZ3BSQ+pi
ZX7xivuJ3HoBTPtKWJz9hg==
`protect END_PROTECTED
