`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46hOcKrGa7pL+3HdJMQ0ybVoEmwL1oXvLzxZz/vgII+v
U//OHPMcxBaTCVWL4dJx7Dr7jtJ3bdUwau93m7WUqwcADqUsg3U3ZpARcizTSSBK
HI3UixwqaKgT8ge7bikQDExJ71wDFjwIgYnhz6nyK9o/MiQyGB40oQ7tGoiZ9Ydu
sEbWj8akfVNVBkcUnHFyU1ML/GucIM/iWX19YNFxC0l0WaAlnvyLlAZOh4xyJ/ts
N6wZePvDVHdfF0Q0w8eQYVl7Lk5+HmnbPe5MWNhFZh5mCGGuXnNf2Iyh1YHADe6i
hthi5ln2YuRdjUG1RzWvVdybnq4ETKGnPHqt2WG3+dIi2aqWr3LpPtRWIocpAT8L
WHvvDLsUEytQS/TNWhIuUQ==
`protect END_PROTECTED
