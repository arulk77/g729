`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiK2lyubGP/bVaIiNjCgAcvly6QSUkzIjltUiM3JTTJAZb
Vs58E0CmitWISg0SMLcUTSNUMSqfKiRGeQsGWvfMAoToeDBfsgwqOU7ZzbJxzG3Q
m1xBIgq1w8zGsBM8jcmKWOK/0ylVwu0eH7xLC3lJ4/FuC/rm4dao8GGwC2zINRC9
aEn0P40E8wvOhKMsgmESGg==
`protect END_PROTECTED
