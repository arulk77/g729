`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tb/dmh8r9ndgoP5vFQ5T0cEBpubboOdXd4CvgL3Sl+PYlb4IBquotXYa8nKfOnfO
e2D7zcea7EnyOqpHKmykM+93jTG2nrdqnO7fcCw4dN2yoz0491MBL2laq14aDMIL
WKELI7TuWcSRjSaBYDtJ108YofAzThzRSUTRMIsQfMInz0BrC7vy6kd6AQGF3Bc0
WRXGTHTYUN1xud9kpNwhWU3LBjuohfSumK2KoeOeEuJzRWnbvyo98u4Z0aLds10J
q2hv2E6FcdOegQzb6nfu3yIJraCv98BHiYYgkiZIPsKwASrSrGkquFQLBqrjeVRa
P4vHlAKFN2JRt0+GeKoUoL4RoHwtnmFJ62bz6cWlX3qQS2l4mL7CMbT4BqetwJ2C
DDAwk6hDE0kG4bwNw9hiv+Lg+ii6Rl3sIwxGMAsAQrrEdlCDNzEND8l7/W5MYTpj
uSHbC27EnVw6+Ypo2mrGMo5xPIdfiSjS1u3Ajhi4OQNKMBUuK0empi5CVbVxbPqT
vaVLhTXFnmpIqWcXFlExWsFaPPy8gMv/rQX95amG+4+mLpk+H2ZB8pIxvKQqEzmH
Ds+QZCQb7Ee1fkWMsmMS4kt4WhEMBvyy7BN3VxEwtBt+z35sX8wObbeVWR/1QixV
faR7yfPRTObr7BegLQp3DidTMMJb5hQ30bMySWGUXeA4GzTTCq+DusNpJKcWm3Tv
IfoxJREaGV7pBIrKDg+r482nDwqBDMwS/Jz+gsEUsYFJFtIKZdP3a8Oo4svJIi5P
S73CvsEdrtoHaTXOlP+2Tkq2RVvFjG4L6HITFWsRvtHRdt/DopEeCnT61wSioFIJ
++UH/ExkQ2VGn7hXXmHULSA5uG51t5YoHWk5NDHHkicpleBdfPcdurYtQwtXN/l8
`protect END_PROTECTED
