`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIkWt0im9Z4ZL1CQnR+XqWPyiyD1OJLyt4pqOyKiIKLh
3QYo//I4rQiQ4dPuUbwYkgz9RSOH/+3w0/lXAI46WQfG/LwQAuVa3zt2iccuIzfy
vMrerI9VHk9ozSJrVZdXBEOqGQkoYJ/XkMUXQWlVdc8uhhGV5NlxGvPFOOvDdAgD
Hi3G/tjRF2fLHpN2qHW8Q5hdVvzR43bbYBeYxZiGp1f78I7qbkCHr5usJGEqmiG7
`protect END_PROTECTED
