`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adTl5DkRmQKMFuPQpfm1vX8r+OxrEzeyhkVBx+emsaLE
JZMAzi0I2yfuwQy1xPhm29+ayhxfuBbEreZClfTV1+IuI9fALDLeldLeFBukjw9t
JJkCr2/c01XB+TFbWoOPEf9Bo/zHi6I0I5ynnXhZOLbhOl31WJ6WrepGQ5gNv3r2
OFT2nAl9yJxozLZjNgb7Q5ObcIPeLMCmoABg6fbXBRMcCK4OtN8rCGLR3b87HY4I
ev9mEmroiG1awRlWRG5VZq8QYOJzge5lUgCQDrsK7kXMFQFcRZvMNKuZon832aZw
63zSlyTaZhf+2xR/eTGJgA29jLKU8OuFq49J8jzFs8cNSx0zMrpZu4x2bSDyOyjY
BR6EDIKi+8D5JiFu920m5iJ1ySGwz4YTfO2AMloDjUguK9HBIkqpTmeuIId8TVxC
iL/04kV6tkapGcExbsC1CkCYnWuKReeAcccFjw5pDS+6F4voQSX+hAusx72Dq2Dv
IprgqnPZX934+R+pblWX7Q4OqoN0iowv7OIW36vU1Ucl9geoqpjmfY+KRJV+Yd3R
QOMapXRtNIXsyZYPeOhOgX7cGk6CNXN7Tkp0U9wXVs+cfxIGE0fQyypRJM1ya0wf
dIO2QG40bH7soxrmTCDpKC7PXqQV/t8GVo59CMHHuItFcPDgNkBvHLpxzx1n7A1M
bjuF2k6En1nvOGYuutrdBTkcn0ETe2wS1jlvcYxRFPJuZc+CE7bVEj8+X0SXMdn5
ti/tBYClSi46MhMKRbzDvnIQQ2MGwASTjrzN+QpDMJ1pBi7YufDYaIwdPP1cgQvR
/cmsjC+W3Vd5f+yvOO0yaqHklJNR6r8tJAnPBxVZvuHnvN4qWmJsS3oZyGsStZ7W
42HEBrdnJZ+KOj9gA+QpgmYoz+IoUmk1rZpBen4HZ0qglbGWX5eaJJyPSVYau7NW
NM2u0fli3lcazgCQo8sB5mszp4i/qIemXJsd7k0TdYb68e9LB/wWjpM7AW3XCFoQ
5jDlZKw0cicZetBcsmbCfTGpzu5m5fnw7V4/2hQV01c=
`protect END_PROTECTED
