`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkdMIEVrAbN+LNWXt/+CPL/vtQOCVDYE7O3gGdO6G4m7j
wr/y9IaHNZBIQJulH8BNEp2EERNyLOW2rRPNfA8d3HX4aiz81pYSefy/DjhCoSTk
Dn07ZDaFNQqELTA7z5GcTw2qGx5xRdZ41j8AEnxptmDaLE1gRKcW+gDRduvyub1C
L5zImlsesUwy1NUoRZaREJXSK7r/BLMCe0iV0297jNjwpO/i4NN6m61UBTNL/9yS
mr2XbVgnoQBwXNrPSeJMHprcx+4SHRrC3Vnhfsg74ufbGtWfw6gUUgZGgv6PuYu4
T+ox2VxFu+z94NcowVV2oj4u4JLZytN4MoWbN58+IzGLbVT1UktVH+3eM6IRPPYL
69hpkvwVU+LhWLb3lkiNCsMnandpjcldmoixwnAOGVS0//CgUpL9urK+uZ1BsKd5
d1dh2hj+MK60SY3LoaujLCBWFooLvFE2VJMKVcUxdMHsFhv+Xlq5l/KjB55UGQmx
`protect END_PROTECTED
