`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bkQRH75nqJjYKa9DzWuQsR8AUbax8k7N46qPws+GvlifdkwJgUvpVWSni18xWBnd
g7ZpVg+rakx8xGlzdxXZE1lpe8l5bOAJSSRhr2lIyumzOiEbZS2/jryQM0i2VF57
l2CmYs7zQmGYv10yMuvgJSHYpASdg6fzKRtuD0CqilMsXr1ZLy0DKd94lBWtK550
xE0ilwMtbw/cJ0QF8hEbZWpSf9Pe4Eyuh0BKDm2NFKbHn44wnuucccdMVmlvBHqe
26s4vSYQ0HBWfO29mnlBT0AwyfgZKvZ5h0r72CJ8JbbXan3f+0rHTg7IdxP6Aqo5
Pzalui9DRixgPL2NvMakQ+LVLUt+XWG5iBbGJco9AiU=
`protect END_PROTECTED
