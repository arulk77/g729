`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
uIbczpsm75wWH2aiRiy8laONt5NVsgAPJuXIxTkz/BIDMFePICm5578PTpHYVDD/
0vnjFKj3GjEA+V/umIQTGivuq0BVia1Ntj+YM3+zqrLrsOg4Pky6dtzvcFAG/xjF
oBpZ59liYZWrZXk3C5CaPYde6r0JeNjB7bKJJQfyXxwxnMEVhij8Iu7NYIYaIvED
s/3RB36ONxbhUpQQMglLeRsoYblvNmQUx1F5DD2m5G7CuCchVPwJYMJqC1NB8RL5
0iG7SMeOFWkztik8SekFEjLUPIvTSWMXkvsLl5QffM9JN4CoKUEJ/nPoVeztSu4m
fHQSGbmT0Ar3hkMh/SKE3SubfWz6DkYEdlX5y/6uPFKAcfGmhdI9Yv//ICIm94bO
PYS2wp0r38u9BmVhFaTv+ogTYDgkHOIcQY32qzcwNiJFsQ0UjMX/WcW7SbhKva0F
9f2wBII2RldwbEiim2OKZZeN8iIz75AoFiUaaIiMpvqFu0dscGcvWyDTzZWdj8pj
1sGr8lNJ0FK5tLYBIpXYGcxrenO5DCSgxVPQw5pbDuhq+L1vKOUx6d6o91VOsM7K
lK1TGlC+T60w7BjMB300n5vtJ+suHHBF0DpnM67Pl6wqGPLCn0iLrULAfT4KRwAO
axV+Drj00TR73vNuWWvdXsvWmEQUcSx7rZ3Pbs6Ov8ym4BsiF+mGDq4ehXj20ZGk
`protect END_PROTECTED
