`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEzkv3aiCGuW1Ug7a26hvcak2ab670CMOmyPhsnqadbM
inN9vrS+1YOd8CH8EsJBVVPqImkROWbG/X5N5LuCkHZRhy3JKRKXmVAhaYWXVrep
aYz7Ws7KVC+xOREmG42Yfq9XiwRQ2ecDL7HJ7SogG1nWC10jT0lXAzjIBDvstO08
yn8Fd9miS2D0H1AIcmwd1rvopZaa+2/BTXl91nLI2ThJmUv5YY8l+3I/tuuzWBhq
ToCHhlRFv3EKVVm0B9GqTV+0e4i+Ivp+ifRSF1BzCZRAqz5SsUFdXLLuoIgehIOD
d5x/99nENPpfy93qFzkH6t6D3p89c+Gr+WnDF3ntfM0xnk/8sTnlBHVDe2tA3aNy
`protect END_PROTECTED
