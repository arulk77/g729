`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNlxwIZ4loMsiJqtaEGqWT2K87QT3AJUnojAFHwVOba8
xtt+BFh1eCkif4wdYHCi4GIGrkiHXRrkcLOOAd8mlehaiLo4eff/7rXhfBmqx4j9
99TNSloVGzW1B//1U3A6V6dE7hbsN3xpEEs+6ScxyJO4tPkwInfuI+pkl8HnYWgF
Tiuv5PaWdjoSMDpME3ylMs8MlxLZRUF7HDcofSWfx53bmExwLM9OxUeUgUMFi9g2
EADQ/bmydjLCtqQv2lIdC8CYx19N6+CQ4poQDjY1l/7gx/2dME9cgt+++R6Qyey8
Q9BDeTBw9ELRSr/3gGFie2A0KhOmrXsVqb+aYcvwZkKufKXOMRxn1yXe8nlfoCQe
xsNgd5yScf58lxeD15Bi0/YzeqMR3J7DLXCh9iKHNqj0BcRVS1FFA9homEmVeX3g
vFv+1KPkx9y6WoNO7SKWNZKtPGTa3qsqPixc39nKaVUyXjjcBhm6+Tu5oSUj2D85
`protect END_PROTECTED
