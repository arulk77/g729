`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42czoetwAHzhzzJxQf0bBV82Rqnibwg1a7s9BzuGvLaw
N9F8OYvxh2vKAk+e8drgvk8IsR/gehh42MIa1hPnUSl3otnbbBlVl0pUN/HPFROF
bOhy14DXO8+GYPnv+jEWf25DmxutEJfSI1DRzvIQpAi4chyjj+++wP5lyb6JHtNJ
ujdtYFGK8d914eZUS0uXUipoBXNPxQojne99fMRTE9o=
`protect END_PROTECTED
