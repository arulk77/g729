`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QxXGoZtoCW1pbBOsn4vcEKRbL07wmJ/+jCsVfpwrTxzFyz/iIUCW56rXSI0kRsfZ
qZrLAiQpMRUfK1P1Qt+LdE5xrsojId7PnRSsW01bHuNNrK1T/bHRfDiSysCl4UW8
pnpOF7zkN2JWnJ7RFz133EdE297Om3/cuSEhaz/RnPy+KuWjmTKl2bev7hQBjkMW
p2vq78aJImH5y1B1iipULmqFQx5zLJqzmMF3U8pk2/o=
`protect END_PROTECTED
