`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
w1l/e+WrhRNDzXKLn28YxL0KEiZeHqwbPzQ11vpJ1Gb1FI0SNPzu3ux8JuUANfAs
T2bIEsMaJTuho8QvVbzR0av0yoBVfl4QGGvn6riD7PiqCVAc/VX/EvG7s7QKUWYA
5VU5MstR0ZuqsHyYJJF96chDPHb+Z7/p+zAtbcaKNQ/WQQqcGVYSD62yS/e9Dxqr
oFODkACj/73f5W8m62DxTKW1+PBlYHLGWsjdXYuVfOdwcdUfoNmagmJjifsYCnx7
kf06IJFU0bsUz3v5Lh8A7TBWp+DT1UEEw5h7qf749jXgs5Kb8Rq5Xi2aAIAqitdj
FVbCQJjJgDH9s8N2vepL1012mHcsXMFCA5vlAC41Kmymk+cqcAg4cZen8G42N8Xv
KRa3cjUEnRy0oHb9fYQvgwBzP05rORtINiE9W9I27XxL6FJ/B5Jz4jkXyWlpAsV2
7ns+BkV7tT/L5H0I1NPbjXRD6z3pf6P9K7sCvpAjyn5SPeBqJv+qcOEAjywY5y0v
meYK+01We1bgn88gTyL1fN3osiMdCfP2/AugoefAFG1SVZO9TQVqL5yXVFLWepl/
we9uWLAGBZle/LMoLy1tKri1LAfXXrdB7bpFheUMRuvq7E3OAwRwpQeJlIs/9YMp
g/kgAbsTzegjM3beimakQeY/vOCha6xx8cmusVFlNy4yBep8f30s9nfU4t/oqZ+N
sM1vdbAZLNUtqOw/Ti3XkUZC2wKtZ22MSusamdxa3OOGfKGaze1YWRz5zD2V7ihq
JU2O/WoSrgBC6W/VKWbjABQD8W8+kSsQCdS49nDdnaGjMDI3cF3G9MGZXEvv9vGC
d2XoYWorxcL4HhXzrvFH9f/h6RpQZB+/j5/i3GB8DWnZhHjPoAHxO3K7VuZJHPrQ
O5XclPCFxgviiWgQEVPqZrnglZlxGOEY5lvmL56AXdsAhFmledvcRlIlIVHvf+vr
h+mu57u3ZD+xAUJAXkVRvLTrHzFuQ+EWB1Gn4ypv+IP+ATsB8Hbf9Bk2bma8SjmC
xXEJqTWx8NqNzLcNjbpLgy6H/Kb08nJe53IY57WJnsrUvUX/Hi8Fe7sBXXH91zFU
Pk648GiXAp0gZsiBYE3T+YW6BWQaTZBPH5jr0tEO2+xcMzDUgvusf9HvrDHwoIfs
TOZEeOj93tb5taqTeaFMHRbGm8kxZpvGYVlGxQeY4fCwmGkq47D5i89SGPkFn6Zb
7/MZHrNq98WATNA9s4AjLzdqjG/tq/yE88Z6g9YoigWmnCxKZFWiqXOToyHRM7UP
0nGjEVgcj0VC5oDp2SPH3Y9vU8Ok63it2v21P84wPRwL7kDdWwlg1sK5eJlCX1tl
FC7gRj7RKIkMYtNQyUh+7F5T1+RJDM/6pj/DZm1FoYsWTkvB7bdOBBi8sr2kNgUr
tl8fAy+ouh68gOli2Sk4VlinDpXekgvuIsde0VNh34VOwNbQDxS/wZJOVrKVh6KI
npDB7PkXM2Z7Wl2sww9fzDFW1SI/XgM6xPrNXcYMNTSJvWNx7xNMF0LNNkEuZpWo
DvJiyU9Y6fagdEZVcHUOpfCetlCB2ifEns4FMd+2MK/WLr5XRVG9XB/AP5xXgroa
A6WAP6dtfLlFifd75bk5DtCByJZvvd45Md19J7WNXFZZ2A0XCrevnsgTmc2C8f1Z
+h4TB/5hCXpjurAwgmLiKCgHXSuDGgrn+oXDPeOEKsdaI1N9YbUmN7slsnzQscZM
g+2Byr76NVjVTTqedajaNzQXqet1DGN6cMmSede932QGhEfzhwLepjc6un6nYUUo
VrptEcJquOODeAAqP7ZjjOVVGJ//SJW4lsr6Gm210EEFp2NPB5lgBVUZ5JqIY5b2
7DODjZNyUMNJHCEWAPNFO9XderLZWa/btOEwcxETqqKta4zjlRhYHHY1cPTOJfhD
RgswsWu2KEp+4wunGMaKAHZOZJNCtNmz8zQNeqcJK8vP4kyDzmzSwW3EF15O0v1b
EH9JPJ5MDEQCOQRY36UwNnauoUZoln8aUymqTAlJMWy8tcBJ3WtBezztDNv6/twt
oXBw+FvS8jnhYeQWk2ptV9DnZkx3SPStOUTaMgJqWB0RjBW1NLqTcYiyqJVqoJ4O
fR4DGR7NK9PlYcBvSbie3iTvFTOIAKIh4+92F7ya9j8UnpyBAEXPZftwGmBQipbP
9ZT94T44cQsciReL8lPbIgCM3ndU0hms2HpPEw8gbygDqIKGuzIjwRTae4aKlkX8
CjpMONi2i8EqWTPx9oTXe5g1Ej/IeW2c0uZ6m0ykmxHWBxyPr9v7q+fMfaCIQApT
eV4S30BhFdF3GBi+VBkVVObDDdIIcGlp2PsRw9NuANar3vm/rfNNUPsfCpA6fzDF
N8BowENuxK0+ts9qR9wMy/Ccz7rbWQChIOzweVOQmm/PPK3XcFn4893fcO285x3a
TymL2J/BXndtmJ4K8ypz5MqGbK+NnGxXqIwrs3yu9bGoGQLovGEV+jJMVwSdb3PZ
Kx7rcRsgtxQqemyOPG1AVzim4tt87t4TEvGQbAMLLvhl9wdSwADxho6c51zBo7Z+
1UaVDk2VtPKc5fblzWmcwPm1k4BDUFfeOUydqlxn4EphC3b3hrqjdWeW2pXz2YMp
tNaf4NAvHrxHpRmIQ9J78/AGNFOvHkkcMSyVnpSEXtsv4KTSgcgZgi0v6I/c9K1H
SeX6wyOroNtRxXRl6j7u6n3C26Cv6VcA4yi3cMTw1wX7ylkwOZav58DBq/gBm00T
/MGvtynp133sRzTthi8UzB7TZdn2K/rwK/rLOzyoNM9vkYE961gXwrySYAvyXvDE
HVDcjk1TFA6w8fFC7uHLb0bBC4D9D49nzm1jk+pb9l/Q6XoLXdj7du0cL+1WDRpz
zXM+LscbB6rNcvMe3x8AyUhTUsKElsHAZDTsidD1v+mXCRsxKK8BGBBwsDV6guLB
GegaVMQh/012L5lifvgof72LEfi+UC8TI7flWeQspBz9xqksZr/3CAJPNAbHG4jO
uO5hgJR2qZLsvrx/f3OVNecynRjvFj4oimi0nHIGSUV/12gHvukRBYEHMf92+Kca
Vv2wTVLfYB+xxBpNfqz7XhlGbLICykGP4dAA9uJb59pnl4gPm5JDMQhQX2zlWMtg
iTaQdnDb40vIk+caSEQVs10kQztBLmpGloGlYKG6u5rH8u7qd8YxKN8ffAjdncnS
wKQU/clw9gMcxSEK7O7RcGt362DQ+dICKUcZabxh+VfO4G8At2OX9atpbVe1yhs6
wmipANxWtwQ8e4UZ6dJj0A433ZEuCH3gc6J+TwpvyLfNkeCnsMlJGj+xg0u6ao7+
dJmUZOMAJHx/w4cFFX7Cs7Kzwk0sALqLHg2iBwzz0kIQKvrrz+GX4YPEquIVzK+O
DN5cgpbq8FRL2tvkesLRypg95ZTcJh1hLzf9UXayZ7Et8u+8+kvc18Xa0lZpjkBb
yq+fqKHNfoUIPRDAO1SHOsS3X0Vas/OFX3WWNTIchT7vAANfG9GyItzgJsfUUOqj
bv2iauS5zJBOHDxlWVmxrSvNjPE5nWPh4IY4vudxiDrRh+WtstVjAuGDucOnzPAd
N2THMuB6OA8dlQebYUZOhXbXVENePMhB2y/Zzx1AFI0BjrzPmnVY6iEb/dTJoNTZ
pcW13t3ii48fpMuOujP9nrZhuf+5dgFtpgfQkDCijCDRys9rO6W220fegDlJnsg+
vAT0EKqa2/e32dLLz771unudM6MgTYiJ8zgSHEcCJ5wOsiLxOlQYMN20jsBv9o5T
u4ly0mgzD0zD73j/FcRmi8TsTc6mm9ys4+EDJdgmJl+evWG/L6osWAJlbxvP8Tte
8opa6v+DlINPt8hGNOYdnxT1iM8yWrY19uqFtPFLxOZ8oeYIRt75wIhMLfpUvBre
XRQRrrzGRp5JcX+7jJpsiVC0NsJ9zwg0n28sq3wcLn8+dNpJ4Fz8nFfeJeHPuzvm
52P+H6VCPZpd5zbqQ5BzZEiQ9hVxNfgRdEgN2gIBJOO9YXzrYnPEKeXvj3qAQV4c
oLFit3MNlJU88MQHPNcT/u8+I6eFkd2lutACFerHW2A21IDFFG5cWZ6qUtD/dfvh
Cn5yzxBKvlb/lF0C2jIW6qOQ7iACvjax1B+liqJza75SJaV9JP1aIQmUee5/+SWU
W3GPyeOTG1x0kS+jwqL6ETXAr7VkOAs5kDslHTtmJJUU3Wte7f60SnFlPOCqgG0X
nC6Jz3V0W5Edtl/B0jCnFcFvMgohsKAKmOn3+hcw9S4dub2UJOeu0qcmOzWnKkDF
tfZhHbiLpu63bfnCphO2uo6Ud4OBf5Sw2N0uqCT+ffLN3qSTJ//j634/8tzZ8slD
sSeAtsmI+rgJGukWSDfiAK/HD1BxSaRtNUOtS3iGyYxTcbqfOIXQHfbfHb0WhPcx
42Rrd+91Jgunv1jDbAXDNk6zLuj4CrM5Ik8GY2/oKiia7PWyywWDynyZf8wvOcKN
meaVOVjBRCogi2arsnCcjcWv97rVOXlPo1zJouyNynvrj85zCVlyuy/J7OPwpHB/
X5Vv5R7jweebne1SH1J2+WueBXZVxZI7HKbaxUbB2hRflc0qfmpVtkujrh8L06Ss
WpU06dAWkrrAexXjO9lmehaON49t8lwIrg3iaUZCmQur0IX3c26KePbcOYvy/fSk
mD1iXWfIq0OItcEMyM1EGsPfyrBAbJPiioW9m1AXJleQwVRLzddRULwf/OoHn+Z+
wcBneZ1ZymVfZAfeKB9724VqZJUgk8y7tAG16CZbJnWfc9nUbjsz+ePVDBwp+9cC
A5++IUbrXm2wCIL/9GILrUW89J6ldbWlu+19CILvriOKXMuaECtzjrBwpk0XFbi3
QZfv9KkFEFj4V2FSTwMG/SkOv+fSa5YtC4ivFY79iviG4EB33+3UrM4QU/VJA3Ji
hMEyo+EjXqg/iC+1JPztahGJvNh5uW3tmLSxoCiTPD/9gFt3Mw3BYtym5GTrD2y5
Kq4ic2Z/JSnDxHioYfdais+nA/rLCLkYKmrOKh1lJ38TqkzMfSD48GHW6o960OWC
XDDnhjRRp03R2BTS9tRB1uqKo7bbq1vabi6VEQxYCUopNF92qFMwDJkKQd6X1IOG
z9RM+57DgnhqXBt60kKfoYAm3u+AGAoO0SS9a00MdrnDCZx22xj1YZNVxkZNx3/X
iAqLjO5pRE9DKnQDOps6kspABJxGoS5OxbbTcZ6Dmg01+10iErRdYRFcT1lfF1Jm
P7z7sBGTM5yb+tFL9eMMMgQpmQxSywXtA/JJDoiVT9ibftxAbIqPLSHwXp75tfB0
Kx2k2l33XWmfVYDHEmyzQoi+h4MeozSzXap463okSCAN8VW6EYeFiv/f6v6qnJBH
TZiGeTrksqKH3p/cIbgDzgqxKpIvQGz44XZPF9KkJ0bb4OEqqDgOjdpXguMvFW31
dewRGvfNS7MRVMyHvE/iZTBPeaKPa0bCLOWkqT/1ONsMYyT/edEGu+38ivMmdT3Y
9WBd8irtp3wCAuuxSz6iPLz1Q0w4phEJfguTwH5qnuGx+Me8yaGkte7UnrorTc1P
nfG61FDjDiYZqghuDh+w7tfr1W53Wm83gdr4c74G4V7D/RUTZsyhpsoCtcJbF3jC
EwRJ8JuCMhLC/krim3ZJMj6YpaYJhWgolhH1baY/Gf4WRmJwpxvZza+z7yz23Zvj
hyMWIWDUt65S6OGIXmAYZOgINzXJQgmO54Gm8tAIFhCrck8ZNe/KiQjzil99SNvX
M4SdoZcNU0tA3LYDlMXJ8Gj4WO0KNiHhl2ao/g8+4tMtuF3GAwo5cTfpi7Mu9HKO
6bmEbgj/AF/201j9x4KunpgCGJeUPwycr5liQ7sVHvoaRhTmFPuhZW8pHvS7armO
QmM3MuXes6VEFXefQb4Gqo+lVbmqozbarFZFB2pqdEm7hJY6qdQFYXteG8oFsRoa
cIE37pWJpNTE6kkrQd9mRWRMEDx5iPOm/DSF6xdw7pAXRb4pY9snPnQJSQqNTTyG
euOu47F+FpeAxJQ9dXyUX6ad8tfmhr3a5xHInnWwS/sGD7Vrdjhd46xitIPhZ656
iL0o6TKtyMvXdGKT2hHRWOCrwakgXHfPNadHitu2nxx9Jkw0UpK0TA9zaXhhoMQ+
P61fcoLuB2AUZwYDVhwUU8UX06NenwF6kWBvjpC6tw2KbqPs97MHVU4ZEh3KCXi9
IivRq9RHgyF6qjerlX6DEY0vDFPNWMEey202pamf08byw2LAE6RLZhPsbWX6FVQk
DV+4p+6tNEdr61sfZ3hgqq+GxIOBn4Gs6zcnqeYO/SNTnU3+p3AO+r7KelEIRLJN
bDuihG/b1+vJMZSjSXshO+RF5j850+jWSd3UREQb4wm1nV7cW6RzsK7vXG41cLG6
YkC0eaL5agfo9n+qSyLRYtEDhjJFoPENQbAfpdefQdXCAt8foH5II1yLavfcN6qT
s8WFQ8Nh14qQgfqmGyskNMm2aSFKCrkf2BEvaOMJf+9+VlEhzx8PZljMNNfQ7BAv
7Rti4mrXnGWHVHaFNy6HA65yLkqys+MhnO1+n80GAOYAGCFqImf5lXzBD3+snmOV
X3WU9Oygcfw2DUhG4MtwtBzVJFZyZFnUsxKlEohKzBBSiflrinN5WOgjdK7O0/7l
wu3Y1xA+2uHNyCoFQEep5qc6zbCUYV4UKxdTEzYJKNrdV/XggN5aMromXX+3s/zx
AZDgQGGA2R7QtaqExUSfxWmuvvVZsZXqlEpkmKYY3LldABe003Holws0GoLX5Fgg
iim0PztCiXp+9sEKiDKr989upD8Cqa1EqOxcGB3egWjMg1rv09FMYZHKGhwAXkWi
Fgt/Jzi91hLjCWTOCYpxsbQ9q4oL7ePc4Is5QQqNsZx0WfRPuADENzCr8ElPAyVI
0TQ8XgVl916M7sQ3eTb1jrkM30AMwx9wDW6NoiCSA4Lk7loujpqR1ScGoPM6OILY
j8fQ4fMVqdwacqc24ToMWpF43NcFewtNRzYVcAsJ9Cw4CnW+wIjtuagA8fFHxSNf
AE4e7W/iEfdx05+oWAbAdk7MdNUHijBcCynJDoClKB2YgnBS+h+bUm6dU34STFQs
IFvJjzjL8fLqQqkmk9SdaZDdheAhVgybqA4abR1ArfEs8KMKKQTCPruS6EpMiUgN
Bq+ieBm0EB2L+pYds2VEKqOLqFl8wlOiB/j9ryhvo7jRK9w00U8ClVT4RnnyfKaN
Vh0G5keZlI+K97X8QwFfg++nZi+C7Lp7SFfrCcHnwRxAn8tpCqthpddEC9Yf5VPR
lDOj1XZABaJd5nAhVcpYtlRNLGYzD072G25QpT9w6Ib/9jpFtDCjQMG2+nco45OM
QxbOoA4qBwzdiOuEdvL2pXxRtxQS5cwVOHwyPzpqFAlONnUn7dzRKvTpsY3bMrdg
482q8tZC4N+zi9StGPc1bOJT/14WOk1oYTD03WHh/zRgck1evh9HChA05o4ebmiW
ONUX+v/jrz1TU5xefjgqmlqaHl8ZU/2HdiuFb468vEvNRsrohKONyeYaBXu02CcY
kYdUPGJH5NdJAkPyo+Q5Z2m9KucaLCKpevnzeLgvl+QOTU+7HHh4mhBYVfc/bm7s
ffF5mPbdmT9VTDw/dZl1jhkbPFmIRx0GZhiiDtlWDnFPdETZBPl6HW1kwI+7Qkrg
ovMER5sGkBo+rIjlR7w0AbhPKC9Y+CiRVxhA6FT5RF4tt683P6pSofM3fD+dA2lh
WaGJpeXb/S2sDoRNDxMnkndEC/uLGkLAQYLMw4h6QVU2QmHedND5XOF/EQmhmtc9
kZdt86XYcubN6zaebxp3C9BD7apJKolSJplAwjB3EczuMzL8wN5PzSV7ySBtUQ05
faA2a2MaX9OVv7jIg5GP4g8u6P+hbSht/HzHA7wLHSQCVEr8gDRZQTTMyisFDqNh
tuJ0/vF9NXafRRaAq89ekJ2dpkbjsA+q2UAVnaZA3sEIk27Ob6D6RV4g/TeTrwoB
MsWuAwAmR2/qTvaqUW5aI1HAINRvZBwo5TkH6KZxeUCxzc7VjfIB0IHZXIUWDf4P
j+iqzQI3sMo1pv1JwYM2kCPkAa8uMBkYoJYupbzjfjbvdVQ0zCoRYBad1PEZCaX3
RuiZ+ga/8leG2qINfmcPQNPhb1rSKG05YDirCq+0VXyeYoOY9Bnd8NkcZhJYfN7X
Sk05VP9MWGpuJ7XMieIqOoPV6+izhIhplQX1A63fJjfuTKI7GcAorn0M8ywVBriE
8y0FJ/e8hQEHUpnuN0l+bcdT8UYfGbfaXN05UF3brXn50qXf/bdIQJw/emmKDoSY
jRTCBJXG0gwzSx6Gj+31QDJYcZIPoiUNTUPPN8eq3vUebG1t5qjsFF2oRNHCBtgY
AGPYX41N+7wv1ViNGpeS4IDv7+keMuB7QnyzDU1mbjGC4+8m7mOHgu8mxAJOvhab
3PnSBT99VoxXN+ygxft2y5IS6d0VN5IXayP6A4VSOb+QRVlMyEm1ni5fIxSwvXs0
usbeg4tlh8vpYmZBj9ikAMFGI/UNtcLs0h9rmD1DahZPyJGNi+yz4RAuhT0OM7b1
ZlfXl/PTIaDbf/+W3Xq2hOlBbVFO37pbYmBqTyfuCkFTPIDIqY8aZoqllj9sxVy3
zfiejjMOnnAKcdGfa01O9FUlsS3H1AqPh3qIVefH8NqyHKPWhnxIDH/ShkvSKkmf
Y6+Z6nW60FADRYETZBFkA4iu5+41MCNszYTXJV5gxxBsIc5jicL9yPpQsqF2yp5/
EFiEvIBjb/HEyUnHwNyMx+fKVqNPiPR8vZ5NjSf4jz2FKAZbRvEgoRUTUlq2ix23
nmb97P3xc9m50gl4SnjPQNbxoUaiPwmDoqdoTEo6wS6uIOfTu62NaEbxv7oZst/S
os7IbOhq4p6usyA1CXeWx5C3+kEqcp4flQhOh7W6TC60OtynZoz9BOGDHXTDtE6P
noxBqLuhOllEzxF1SkpQQK+GToqlFp50vDVdC3yITFvmQMW+lIioe47o03m5x6oa
JHtkYk03dlPTn37l+ULM/Nmic1MPj5oCLdz6VE0FUX7rXrOVTwYJ3wiWGSFP3SU3
OIWpCppyVYBgkLKV1It2fBq6YxN/UfMFIPjEFrHQdzttR/sGA2rO263sle6WcwEZ
XEvy/7wqnsGjRGElKVF4c2I3xcPH9DEQVUVoPD8dheqrDw5KoCzhNdOR5ZDqrNYg
b8pGXLI9v3riQu3ySFOjBoc2tGoGmTCK3FbJaCHryD1BD3mtBUBNIDMKnqNQm7Jy
7ZmepDRhNxme3MmuEC3v0bzXbqqEK2AVwg5phQvx0L9vesrpwAtK9nB8n36bpqYC
rRQKPx9air9UBurk1UampZsOjaXC9xmc4AsYMgXQ5+qovIMQctl4lpfQImHvOrO2
MtQ3PC7wN3SLQHN4tV2xGb/gtyTBQCiaULB0Ts4gXmnng5+tYoNC1p2DbMVLTKDr
BKKCDjLerBMlcmFkKho/VHKVg4w+LBTlFBCbjQwxaZaIxQgepCGhLM19ZsGCtPUw
Fq/hIqyR9CnlQUB7bmM7pOuX1XP5YqQKT7qMKyQB52FXuHdzYQG875OmKLZVG5hk
2lRKKcBFwVdKwlmlcZeZjZ5mdEfm2l4GEwkCw1YFVcLtWV21P9R5bl5StOfc4QM8
VLtPlto92e1Rj454XnwOCuppaQj36agll6BtSDfBo0EFq+FWnaunmJQvZ2o/X+WR
40J0Egd0NVwMgxke+noMceBNj7EV35BF6Gf9q7tX1JL3BmHDBwHDWcyXXka0b00C
Sg3B7PvyQmtnwCOeclqZI2Mv1JrL+IksqA7KXxh+tzFL45conuk0bFP1dwGyw7ZL
sPG4AADNNlAxdB/SWc1lAzw91SczywJcTrGI4JaeMhAdw3aS7RWtIl3oWnqnJ0iJ
HgCL68TLQHtaE3HQboSyh7uio+pw/hHCA6NBYYLKN742uR6xbA2u47Nqlj12rai9
wMISLd6jyfd9GgkgD6Fyjnc1NNinLpwqxFqZxb1QVKgHCbq6nQgPGbIjq0hUOlTD
4f0XlZMLrKO68dAzuNIimymclkmHSfQmqGaAhLplolsZgv6JpcNJXir/Tcfow9Z7
NPAdVx2qSRFdCFD7bwnlgCp0ngH/PYWcb/ik0nNpC/4uiJmBmO1MOjKeH2dZfN/Z
esJrW/XHB/Oi5KA03L8slRnPSD1+mrwqvXmk1biD+y5Zjz2Bl6vhnaY6GTST+9/w
+uo1oV+X/5HwBIO53pK8QzeuPHMULFPrlIEN2vxh39asGr1fyTzx4bd63NGl0KdB
bY71mmwcJZ9ma4ZyRJMHOjbAHPvkQ/MHrUdvjH5BQkKnjDm9MtIJzMOGYeyNrRgv
qTbQstzfQF6uu4VYw4BAnr7V33aoDfkNjddqojb7H5HdkmOGMXCBl8Ofakzvmxau
qAmVNUILjHONBgTjV7OnNgHhN9vTmLGUkqon3gM6QAoDA4usA4dR4jM0QsmhK5MN
v5eebGvNw53HFwbLFXUJ20gs/cSiqCq/uzKK5SitW4IaZX99b3mCPl/Nps0wCcHO
LYYcudHQImOTAxH2lYqkqgAUbXNI/JjbpH4lursRSxGw2UeUsSrkxJxYt/+Y6XSK
DpAAvNIigUEBTPYAXJ2+G8azXkgB1lsjHf/oZHRToPEKWVxWz1JWepF9+T3BQ8Ed
GNaisAxiAuWCgnJCCTbKgHW7NQ9sAwHwoIGTlLQivGw9VzLZoXmi0QkgWGrIdxRI
RpuLznj+fFKNGvU+UGFhmfvFe0akbOvvjQ2/iNJwmE/bWH4ApRRc4zdEXJ7i4TBh
Oi48u+4ecI/y/Jo8L533kLwB+Q/WbuljPnldYuUmYv2/L6hUAnQXslZBz9EAHsia
PFN5eSlY6x4Roqk2e1hu2JqQjo0aUKWnurp8YsZ/a8qfjib3tPP/MA57E+1/EN6r
0BDwR4jwlyik239BOVWSmY9gnWMfiTGXa5dl8bT2KVv2KegewmRiS1TrObZXMj6J
1MsiM8IIfAIWpIxoOT5YVAD0ED8rsJxBytbKuTOMqbcurieOld7c6TDV7E9I8NbR
W2lvZE6D6YmFoW6vJFmKj04JgMHvTxmwSvafsmMJMaNJ34o4cRp3YQamOFWpMdES
j8q70xDTq+JcZ3qprkQQfFM22UH3ANf7DA2DRfrra/BTCRcIGMC0ZI4yPqGnF6YF
fptU7aUMtdWW7ZHDO55wdY+zafbWipk20phUFoZs3+S68pGpri88KjzWOXDn5c5V
48tlN1B0dVYDxGJVkDlX/5MZkI7kGXd8msxCLhgucmC4jvzL4emlU1aIVcUqplTu
x9OLW4/7DZEk9T1EFDlZ1n8rCkJCNwXnS9S8867M2lKVN052+I+EsV2ielkP+pjJ
YRSg4vtdu+3MQXl8Z5yWkWFuwlR8YYQewLKd2LZFZ8ocEhemAzknOhLOzPTtE/8L
vSJoeS1TS8ilNGVu3J7TSCb/6LvgV3Tn6rIETB1rvFI5hdpbA6lhr0/GF0UnrOj9
bxl7ukN/Hvdy3+VLQy/qNy4kvhzsTTeDmPTDKNFwomZmx2pwfdyE9p4jEZFJZJX7
xclrJbpgHElW0W3v1VsuBAWIhTkgFg2BhLUsJ5EfWr6ObIfHcESbnfnZ0yBZEQrv
STwjcHOBX9r7gK7qboMIf7npgthZJsAy1tP0wIDZdHvZKlJwQ1JOtjGfnZgASKH8
iaKRGQs0KKCKFDfONkRl/VeoKqv83U805jaXE5R9VNqD7MG1hQCQwUpwQYkaunZe
5cwjdPa/pPoOWiyWkVsxb/ki2puz/YwBUv81BhBn4u5gy8uZEYKzUMPXzXgGyFat
DV94Sa0JXzA1nBA8W/qQ3GrCnAyMy3lDgmwYSOs1C6tKfDql8Myo5AEwFPUe4xra
un1Zd8z/XzwiTAb6YfIwWDHlsy9RrpcVOwW8r7AupLD+g+vmXugZIzPMAR7xD2jG
+CSPQ2NLfRNNBfc8YD+oGQPw6oYNXDebHE4b9EhLo7Kvg/fd6ZP6bxTrmsj8SJ4p
UkQQ46cRFBaO713142T2aJnoLqKTdvUFmpdpAmFlcHVHSsbHj64oDucVn2XTUshD
k1vqiHvpfmDMV6+sQjNhgn0Wsav0NcHtZJXs7P3xRqRSA+YogqXY3lwAZSlxAMZX
jqDJvlS+M0HJydOy9ZfmSQIKe7KCTHm5kaRbgAYFVxNwqCkWtFb+2QhqwWY7DR4t
J22Ug8n7y5Bdxe8U1HUhNupOIMjPGDd0QtiFh2mCb7AgiHkNhZYGXUUDzh7EOq26
CVkLHCuTL2L/AcB/AIBYOfFE1Ej69DvCbNmhedpI2iv+RlFDO4cAn+TKv9rHCrbd
GH7qWZ4rDBv4WZdD9kGqLMmlPlQBBFNK8kZxuyO6sAGPgIGm1K+klzaMC0hd0u+z
rOD/L9xdlbRa9bi5i5bYJlZsakQqY1oyjRtWmgDSTfcMfJFGjATBF7emAwvPDGfc
5rcy7afqcpZtbOymMa6Lg+SEONkkry23MInVAVgWbv5QN3PgA+hFDH/xKbRVEAAM
zIH8UJuVpCTbkb956qwnjHakSYNsXOYIS5zX+CbQjsYcZ1XuTYyj1Ef/iqkn7woC
CYgIx1olraP+fun2yWax4uT3oWH15yeiWfHEHJRJ72IcVvRlkkhKlRJCWUhyHsvZ
CbAJOK+7CmOSwp80oVB7MtUsChBrxl3qhD4DSmLRK2IcFoxA/nabyUwqBarA/TCw
F+s7TB8aYL2KvR3lbPbjNj35BcodKEEsRFqsScPG47T7/opA5vsU1DogQJDBSRfR
PHc9/Zohhml9lBRBQlu1g+yzoOaKa2P3/39MF+U94ulWrLZeDrl337npD9ZdelG0
/urJufqa5cCkGEd+/QRgx2LNGFJEZuN9b4JdLl2HbBHJZDAHi9PJO7nkWzNGz220
1xUZbzzHCkaADDKNXCTAKOX9wcHyQmYM9AiBjcu4fhlbGP3bOBmYSiMxTEE2/MAD
oML8L5pWQrFE6sv/jExIoC7q7+MoWb8xzrRkqYavPrY4wJd9ckzdGuhzsv/JM0Sc
fQmxWmb1JiB1nEa3d77obkqENW6EGORHAch3e0ymOmuX/Aw8M/YjhV9lzF5zEgQ4
mVBNLFgS1R80g3lhlkv2f0G5DI8rM8nWHdN9jcgpiJbFjEDcFihPCaNWReKhwZz3
Sf2IrY/ouV9WA0Z3MNScM1ke3EMXXzNExCO2KDO/O/ymsOfhcN2bs7zuJLgZY4SB
cLcZu5ZrXh6Q0VLkXaL7RYNpHTcxylKocGSyzFqBRNbMnVAYOiAiKyMUnXHw/0HT
kPqYz9uh+Hua/+xzs0M1NpQKrTji2j9estdubn6KZCa82XmaNgCO780aFbgM0+un
PCQxnjv1Ail8jV8JV/8KkpnSdEMp4T/hyc2eT1VacZ9JMt9DONSd0qQYCiOPkTq8
bX+tVwbzouqRMYCaygHZLHw5JylqArR9TUEH4AnkVgIz3Bzu3aIqmxYunWNP/e6A
MbilyNnYUa+QfcRqBzD6QsCLq7I+OC8FBExNPpLIBdeKlyiH3uaPNlrqxgXjPxjF
vgl9MT00F7bWcC2Cs1PftU/yGLh0mU0JtRSj2+KjXcQXN+IZGA4VD1je3HK4jVYD
ie/7ScIXpk0r8Bmk4awDf4q2zD+eLXzvNw+JWyXa9FuPvG1v0LOrUuxeAMf9tzjn
Glyzafb759NscmH+E4jqw1IKfbJg6QbbkRK/l5AEXMgrIFYFAoVQs9I3BKR2hu+8
Y5gG5ZF/0kLxIP7Wf6xnXox8aZhDHM+vAhmRPgN2wXxYUTZrX2dRAWiRPvPBO4P8
Qd8lqEM+LtSVAhl+bz4nTwnPwdXL6i3G8ESiN3RW5z6QBq+Q9SLtNvHddPhBT+2U
v4gPqx81OGFDPHu+B5mbp1w6mF0vC7WClL8BUpoZ/1wi1jsqvpaw06zjn+VADVoa
7HYK/zvvtwb0XVScy/AwVvqssXHqX5/RTaeYRyL3h0Tgc+Zl9SLkQqQ6UxNrXt1U
6FFQRsYCxoQedVtrFxWqpXgCpi8PiYNNKVR7UqdFWePCvPMxwheDhlSxazy2XqHD
MJ9JcG5ccinSNcFy5mmi6H0/yidLTc8OlvmrOImfoINTNR9aK8L9JIufkrMzCoHF
hJJCxwkDfn854jLdWPPBiMp7NRSqyRmPqMVsA7PRZzPxr5kYucbXVv6DHhtpWCiV
t9RaFuLPcHSWRyJKDNPSXCNplvPzJCJSVIwvfoXPy+aO1EDTuIAm/+tbDS2vxxXh
fGMbVa+6TKkhNKXSKhH8lg7KrwV/M6sIUMngyc8QddTs2RXCRawEwxFX2lsJzohX
D46IJXkQarZYyT2FzUIvXXloPqrw3jermZ4kppSZk2A+/3lgSEWUioyUBxku+cFE
uVuTiGYkYp1RQ7jHHWzCg1LxRbcFQvBf2ituzRjpA6fybn5Xs06ljtOH+bx473oZ
Y15sIG2/qOtW7zS/fDuoZSlQhWxy1X8VumDzQrcYFLDTzJsP73leYIHhxk7at1pn
nKTEnLi2SHrg+ZVLUupzoySWk30i8UXh93f4mk5tsrVtplvRxNquMqwpDMOf5lnu
+hlvrhQ/yiRw1SuYkbx0bH2D2eViqRrMniCE9Q5u9hVmqOq6ycWFBKAyBhD8wlxs
1H1C17ZdsxmMOnCOhWbIGla/ozUrePTlR4sxqEIjuoMgpo8bxwE2BK2Vf50qJGyR
Bd58YIhDLyIHUyzZpF1OpTIFiCr+xZbn4roIAlKOXX0/Ra/6Mt9z9BNzrL4m8ivG
zPzPQQ/Gra/UYwqPkk/YctCD20A0csuULr9G2wpAGmTDJxiEzl3u3JCbhtv+2PLo
rcEj2PGqrcGqOQizb9A0gBx21bcxzUudomG6Z9GGKZabl9vQE0E2Mkku5egVwfLy
O/1jcQJOj/G6R9bq6/r9HNeTlAi8PkyKlD7PpeyxBZy8EhfoWDd61SO7EPdbuimg
R4kqmqzjmfqnaHEZFrthDz4UGCR5KOeUJl6UIo/pMThOWaqFQAN7kPd1YhBtOF5C
o40MfVXy3njzBYk0HCpl45rC7aV0HmG+2dtGjhXSJ6JckvGHnYXC6ymUqZFxEU1y
v6Bp0PWzTe/CM9o54+y4oQVHD9iYnmkD7IMXT3pPyDPgsUDdosFou6+Hxn7JeXOr
qizMEZ6AsiL7zXyxP7bz5k9C18zGL79m5M9Cmv4J7bKHY14rQ8UZVuKrLJYRnYFq
08EMMV1/ULK7v6LW2uUYmQfhzbRSMlh8Xwn6BbJWfbtA3tx93geJa+zuohbJJV/c
UuhjBBMW2L9ArPvgLAyfonUY5ZISryMVqrKFy1W4A+OG1rzzeHcepfvcdtW3a3PA
2pjJDd0LzmN+QWERHhkpeAw7uSkh2PudaAO4XROdQpyeFQ260Zf4S6oorWWYfnpP
fav3mRObXyL5lYLoxLGo4Id6PRjYnuLBktoYqBUYjEgZGc0QF0+drJvefw9lEtno
l6p29AkmNYdIPPSGQDnwAx1IabQzxg0ik3B2oRzl4dDxKZN1n5H1OLxpkOe1VB0X
PzYrXWa/tvh7Z1UvMDSsKGKUe5qb0fqywzJXHWPU5R3mWN2OTN1GJMnYdUAD97ST
iaSCyB28RVpMcy1F6OnAzPze9b0Y6VE+qsXZd0JxjT1ICn6y5qGG5M7ew2Y+1UqM
anDBy86DyZEW9oCzSacmYDUF6mkUESBnMzlY49gpMdjGDhIUhe8VrBGivL7z6Djz
2h9TI/0/9NpFMkX+pqLEgNlUJPqFKzPbk1OgFtDZ9dlnx32CepgaN5WVJsup2oP9
JY78eCg2GGF8fy6n46EX1MbtxdYoCrrPu3gagOZFIM7uYwK33hD7XX9BmY8t/6fw
XXX5LeCt9A6j63uTTsPHEe9Oc+0DVKV/9aq1w6Gz7jGLGqxlWWwmqbqKvHzjInMx
JZAwszdR6SsqeEM+ZlyGgm1AaR9YiOw5dRwKpfkTCMyQjWQgLFzhMm3xqgR30Avd
NyRxm19JHqLkrVlvExXh/AugEaJ+5M7hg9zSvUMlxpK1BoHA+uUad2lNMFXuVH5a
SumZty3orjapC1qyVcGLH+XNwCPayWL6d16+lj7RGlnZHdQP13i/yuEZFFJMvQla
Tk+93CrSRiWV8i4NW2oDTtWzWsUI1Utn+0q3AcRPM6zDdTWqoEORGIave4mVb4F0
RErHiLddLZCJrLxwCSWvRT920NFKSUVg6tqCrerjDf1ctwGEyCA11Ay1+T7HAquL
h7r2kxtxvcNlTAGuSeIzkdmbbq9UkzolQYjGwky+/RRrx4zBvvAnqlNy50lRcPLM
0JlJ2SlFwvqxZ3zI6oWexucKO4FLp2F1xgjyJB6w9iJAbiPbk05+guGVU7Rz5gHs
2kUk4kBInMQQhHkY6WjEfrzSepd25m1GWxWU3JYbhgDuBJgxdOhdTIMPcqhfcKhw
92gsYjRytoANL+cWwrNFAUerhKvBSQgaHrYhuOP9LSARhvmDyK5wJhKnxOK2w8Yi
/KDznK1louFjfTtTzJcbBO0YMWBKhTAy3zbkB8Y1eO1nmI8rGEwAinB9SgfUXjLe
uOU5W5MzgejnX9yxZ+RDEcaHXxM3EI+DjrI/sJk6zQlhGxbtnD+QI3UA/uzh48hn
Yti8lx0cNFmqpgtW0/Xz5+fWlwd+yKVhgqRWKaaJFUsBXuObe5XeFO5K4OcDwG6q
LEs8D7aEBGupQuYAC0d0v9db93IO8BWw20D/L0DCmX5QxA3+BHkCqTxkmQTQbsnc
NdtANCw3cyoGpY1FEL6PpRhF9TflfoeCpuIMKdCPzRPYYGB8WjbaWT+kREAEryWC
whIH7sxo4QkQePItYBAd1CQ8hHlmSW+wWCgzPlTzhavWaBI8+KBWfM9A/AfaTCOK
B644yada6AM8AjlrqRyZNKWmwGhbIulMLW2oM/bOAE49dUG1N2uJn2RU6A6Jsgwr
4SVGe2WAUZjdSyJBpdvVh5jSscvDo+GbxleM+C+w1sG/ysld0kYfZSeUPw0f/kBe
QR4S/f2P8lmd3P9JK1ozBQodTnTwSZVAmIqseYKzMTR2LJoWAiVaTxESChImpmT0
/rrA2G743GvLoCQltOustwhoKzWcABUJ0F1Gm2j7oLpLi22R7kB0lN1TItSHOX7w
rfdrAHwqp8kCghrfQlRjoyiBpshryUn/NI4Xlul9zPQg7K2eo7PYvmqWHoJsZG89
7aggTvPpRNby6VArPbl72VhAy3dYXIdzmOqyXg2z8M1QyxtWobenY/sGT2IDRS7b
7Iv2oAvTnzz0hw1d4a2c4rMI5TclelhAcYNY4J1oKNVGxkXGw4jOG683mif+Nj3r
SNRiEFHp+GAXDrzdYJmAk1Ul8jw3hm1d7Y2HGawPcUUOagSoFVxjbqWL2uj4TVSv
7Z0mneIrGrSrkWJmkA/P9BS/0DgNKLfZOX3nkIaqfCTxFJTiZwoRoyYWDMPsgOMi
O8oDJa+tBeLMs/m0PAYej6jXbb9KLt5ZBLpDIqsybrvQLrac776kpvBTyhDiaZz2
7oivYlGyVbFbVYdARrcaYq3vW9LOALmml5vy1D/eWgEC11238pnTsNtqmPBW22N/
VcW62nKTrKHjY86GGBB6/U04t1XeLi+84XkFPnfRbqKQVFAHHyyoBnWB0O4TBUoZ
v3tlhMFm6ExfGj1vXy/Q1+Yy1N4U/zWxLZKu6THLy+4oIar3OeYUM5wO29/xhuZX
7doiPAGWKU5OFlQ8eQi+qJ/D8alUsV97NTc3ODpnygUWRfv7iTz0Sp56e4E3ra9J
RMGTaSENP4Azag0YaVGUFAd2SxT3WAaTr2i3VpRXqkrFvQx8AF5i6TIJmti0nYCz
karrS4YmFHVNyaVHMzm391IwjPhKWBs1Rr9R8RPjFoQAKlprnl0/v9SjkWio/GQB
ZRMwXUUh3w2BUig7lWl8EAs+FEV3XJkcb0/KwZfhGKns8TbGnP7Z7Uq0ddCVv+ag
CJlwdJvhmwJBUEvNrx1aVa1dNMKsA9/KxW99tV7Bw1EoI9zxDlGZaM8vp3jiTXb4
rRzBZ3ncPtpzgtzV8T5XnT0Rk3B5dsnFmilk9YIgtKgVAwXQEWzeyPrY2fFBINjz
PejIITh+5XuBXjZE/nYHUDyB9VneSI+UEfhLeJ/fBgxWTXaNYRMkI/Xs4jxBN9c4
RjLQJzJoHb4Hl8PsnUxYbn4kmXtJj//kL5hSGFpEpJgYhL8hwRtepcBztbqZ3GNa
5aZBfXuic/ykHxN5vHkwcfmS+FIxOl5gvEYaiCXQjwSpLp4tpki0wEsBiO+WUmZc
EJ+m1y6RWuHcWQ7b/PhNfrCZPIj4bah/5lIwX6xdBb81dVUi1WfKgg5OYCMWrWqB
XbIWyoD6bnlR7eMhEgh/6DKIVsXqyr4R2w/iTUz0mLUPO8CdA9ohUKWI3jneHhnQ
oolFpHz8rele3JmTYFrQEuEygw9V6c2lyrkMoqxGRH6HRWTPKYj8+kJWDavOMyZx
fpXfNZP2QxDw8dXfkdmKs1CfbD/9mxoJpmfgJk6uX+2EcYngaAdcrgVqNsB4LX8U
sN6yTMhCstxyW6h2ECHv0H1p7ZYO6GAysVUM/pP85/QHQTOk7PA9PbqvvGFEyKXP
6XQ6u9qjG7YViinCvfkYEeHVZwRgLrfG36nKRG8lRqPkyFhBQjnmyPRNFXVJdYjz
goEeVv1F8R1HYW3fDu2noZth+yBt1NDpDrebML8HKivJf/C9Url6CyTF5KI6HEjT
IG3WlwzRoJVVmxIYs+KETWDK9lT8vLf4UbDmJ8nlcT0pGTtCOlcSreZpwQCUJDGw
chqZVmL326kpSky9Vo1i715nZtcNhF2w0M936sGhZqZ0zg2p5bVRdfdXqBZZ/V2A
XH+qQbJyc3/0W/FZjIhiCKEiWPKHKgHwZc8gjwE99R97sTV5oWKUZnzuIwKdE02l
WmERkker0Om7CU3e07MZIowBSd7kShSY8W3bGzLx9ZXEQZaTcP4a3yJauTwqJFYs
Dcn4WWk4vg7pqfFr04QShUFQdQLx5zSRRpodpxtCCHCnjTAnUN0ZjNimHrXKlpoG
WzsWMAfD+b9vD1fglzmMTNmWy86ptAFf6YNF8TVTAHBwkRB0JWDNwOT/Zs4SIu9C
jnSumCIUx2rkAw/NFMvXlLMqV/4zojzVbD4cPeMmfl2dhsQwbeTriQBKlfftD9xx
QnQigewriyx0HlRnszdKvjSYX55LEvjG9u4+/t7QppyWad5ZVrRdbQtC3RnfdzIl
3TfVy5N76Q93ebTX6HX/pWnLrRRRfXu2CWbTmpCYHSRSoAxXTKr3i6+Gfv+IQPCG
yy982zvxDYRH++u2Jo7pg6Qw1JUZgbchxYjiC3y+J9dvma13A3Pe7kHZZGOdmpyl
uspcDyvpOxuGdAmTMmb3zarL0sh1md4MaKN15l4arXct4TTPevN7yASJRBft1Cni
dXyCLAAd7OhUS2CLd9tfdUn7uSpczjtOJKgRlODb8vW/8SiE0xbAstOoY8fP/HRw
a0+Y8tOHr9Zs8L4ZbYDYgpGf3GioW5ieL8yW7Iv1Pj+/jtMAsmvcEAHrzBH9MwvC
JzjK/ZuPAgICbnICArVuVtmFwrFYuvK7qP95BIULq6FNvngSkncGr1WuZxQ+Bxsv
bztKkJU6iUGY2+lx3y1eCCGke3ZQsucoAy1nuw/IvtsJmU8mIbNLcBfOK764Uh8B
x8CT16HB/l3VHypbks6pzyFfd2DSKGnp/94yjY/Ztph/otLJEmplfHqx7L7q698m
nXHZ8dUaBeEqcFxQGPuxUmPi+B5XGaFPS1GoMzrfnngBZ6Vox5HyGRWIHriwHZ5K
qdFlBeozG/PuFOa6aPP3KSF3gXuY1vyksxvp2iMjSRrExT8ZoWqgbClmSmC4jpoH
PwHli1OoLI89KV/Dw6d39e+ndNKRdFvPkKZKlmSgB3nt0LTOF24qPLjiERuVkshC
uRNcNGths8aK3+w10Sk57QDyK4ljBKRAJR+7i1W1gspMqUEdzaKbeOhv7GCBiMgs
pm/5TEatVAVRM3uxMCpym4h8a8lQOlXl+XdZvPvMp6Py3WVXIc2JPtQmryr9k+az
HJLmW4yst1vb2v5SUBOGfho55k2leNb4h3RHHGxhxMcRYmJOHIU78yDIEQ1bsro5
WmyV30OHNMdN2Vbv0k0RsEL3YKmkgAVbtFyVa8IMjNLKX4VK3N6DHTTDIQWQfWSA
idWAzUz7YBvqvOxdM2atGf2/CorCemZAfu1JKXuHuk5dj/jRJ0VWq0WLOVSzHr8U
KcLX2Ej+7hTh+kbIiS8lNPWGcXTsACf7850IH7fVGMbzHfyWV79kC0FrTewtspju
MPPNBTm2T+R4jp5a0yS23LErEljCtrg6OpWKHLHG6BxIosuWMpkvNs8BR1z1ZxT2
hO0ygrDTNa6gJGMgTl+mlcAzL43684Dm0oDYmhsNc9Q6Hv/a3f/EKIhhAGIXwiSd
wUAHJ4FUM6tv6iKtzOQ5R3lHKM5xPnqBIWTyntML9+0BAzZldwaKG/yqaLtgZxqg
VWmGQWMqVSQJ9sE8rIO+8HIvM2u2fhiyfklxLkaAXY87ivC7QvnNurHyavftxsza
okdj6qMZb9joPOOUc+sWcSthKrZ4eXbmQUMj7ugc8gwvP735KaQa99x9tm8SvM6R
wQP5UWqwyKOPBXwNpuSP3K5h+lr7v8R1PC/jg46/CF3BvJXUoymg8HuMOg9OePfi
u2reTtCpm0ttbBB2nfNdBrh8ppeF7Ew+I9aczYV2CaMkkuSBmy6HQDkWIpPvd/1q
uK0hBAaMu6gLwgrVOaBaYa3qhih4tjswfFc4IlJqLcmlsyppD8dg3g9WvZZeKYg+
bZvxl9XKckUwbdYj8v1Iy8hvdsrs0fm7Xy8vdsCrRree2ikWewXB3Y5WVPz2En2n
hM0GlDB50kqY+eYU1eCpGaMu1g4uieWPPyJv9kjIcW4cm/ao8+Z83dstU0JeieOL
h9i8edzyqvmCnojNNZW7wq/NrfgG9090a3WK62vyI5EdF5BHdU6I8UK0br0Uou+T
N6lE2xpcgj1IDjSa3yu89fWvxdZDi68UVYBgzRFktXxfQcA1Bd74x7lc0O+gcjxB
8wMYLWRTtQasjTBhkPf19xGfsunZcSGhGGDZHKS4dtZsBKkFwg0h87cYWUwGFMk8
itIwq5651P313vENIyMie70F1lgAvSAmlj67ykLHiSIarBNs/h+tRqOdDRKbGRNX
zaxnOH0etib6AOmvlCRid1CR8ITDlturqIORnqk5d8X37I6Vn8QdNIsanPibD92v
xk7sC5jhFQEFJsfZLMb0l4m4Zinbwi4JmnXJWVVf5DuHfTORDdWtsnBRy0Jxjrik
3zX3Q6W+/OKD81cpWslOGXFlx/wZUfdLqkNUx6hgnF6svmXN0acX+b7D3le6brGB
OFDMqfgX5ihXrsXWw0arrNH+ya/wCk02F9nFIz6xT/nNXzi2TnoE/oobaHrNn9Em
UKkDSrX9sI8C8XmahyMw0SJ0CqnSgHZdYXiqKyno1mkM3C4UyZqnHJnjogaitmtY
vjY7fmE9pN84b6BlotMxuVz9SFzNlwpiWkkeQrPxvS/51jVPoxu+8Nie6XdaKZuu
TrozpVCaYk3Xuah7YEQc3uo82FvCO5/YKe7f9mmjmiqphyO+xY5us3ID5gIXC/9V
Gs5102/fl9dW/X+PyFI+pfvQQfp3SrHkdsIOSUyhl35yDs7MISNAUB7gKDzJm8GJ
NHOCjZgAOQ8qDBpWr3aTqQiqGqdxrzz8LXFAFXUcQhxwiCw1W7bfnMXs77DFgXUN
q9exCi0xMSS7bjaqZTe/MHkFkG7/lFe8kngSEfa1vTcwhE5piOm0IP6dsylnJtUr
t9Es9fg73Nf2v5iba2cNFj6LcqE9x6IuG5PNthN0jCaE34M17tmg1JZoO2Vv5+aU
HbqDfWDr6LyvdnfQJfhZaXE7I3VjMxukmSs/wtP3MtdgHi5AOjETupNYOCvkzoaa
EbL09WFfVLm+uBuMPLrhMnv3mYRV77zti3yCtaw/mGhsmx8CukfBDde+GJgF3mW0
cBH3rDXSX+A3+nY1NmxzDtUQsLif1k8rAKT3Ob+eI3xujcxR8z/i8MbhrCYhV+B9
g/glARZp2jObhxVfkRC644NoPpuH6ekOdpPVcmdQN1tmJYcexQBytgAIzO6rl+OD
sGqNYDMnS1WVlfXESqTQxedQ38vJziuthF+ceTOOJPU+zYV9Q7y2MImrpOKLk1vj
f7MoWyvX+uXL1T/E1JNqRwiZn+nERbNxQALotcRPw38zxeUYNvlPeMHuim0FaYmF
P6YA+FWtuqcgsFBFkloueX8hY2BLRFu16MYjX1vgqhX5rZ3g3LASDaf0cOXJq5eX
P0tNWKvEeA6hSFuDgpk2KT+M4F18Vi791XdRELFKJRmNpg0VQhlwv5hMKK87FKk4
R3Hey8o84wmUh3/+1faqKFP6r7B5/j1sS8+MguE+Yx2/jW4zgEsGS7vEHAmdkqqR
73+ra8v6B66/J6JubtQBMjghCc0JXzh+iU0Nd7cJ2F+A3ruPrq16Ka8L2Zq1oTLR
/TnZLHkLkVCfw4AdSwZkP1MjX2OJPuJaEHL3SVJp6mzIMSD1iO+YCcxMRCPOnfZ7
UdFRjNOCLrxNeqKbndcZ2wz1Y+9ae68soKVx/CR0T+EyUxKviA3QNI7qP4FtbWkt
v6Nc1dhxIJELqqsGEU9+cCQ2t5I1Hrb+y6O5KwRnoohMmFbIIdVpEFRqiQa8EVoG
ytBEepGgHWmPDNy4eYFAJKHHPmarX3R8cJ27Y1pocropy6koRtflkIERiZTgbujT
VoTCZ+QjZTcK7hQKTkzrS4F+QvQar4qNyBBl9sG9TFSrqIsBJ4LIAJSZtmgD9San
Uk0p7VIf7wtScicyOq5w93IprEHhoMJbnX78HHlO7c1IXiNxRHg5zrYJrjiL/wrA
kzTkCiMuQ3o+XsBNTyVCPuT+X0cc9Jl2vY5NZ6MOZm2TDp4PpPPpDKDx4xoxxuFk
bMPLeuh+WNhdc/miG2lhivcRSGX8fJs2L4VU77LICC+6fi2aEI0a2q8rHT7ldkVX
B/f41yZP96nfAaUVfIlwmhXwiZgk3SnT2xzGDWgm7JL2w69HAAjijIt4PqX5DhNd
ZkDNf0XNjItI9TWq5Y6qDI/XcNAi1F6f1e3a9PY1OsLO9a9m/5+y4hQw8yKY8a4o
BHRaoJIuX5qwMxs8g8lI+nZLE8CfDwSeLkcY4sLEbKPDeSUBmMnQ8zEell8/FS35
tgrciQR8giBksBPxvie2MgEgtXClbHy5iLCfY/kcxDpcf538QUDvHR50EOlPTEa8
z/YRdfcTMz+wei7UvFTSYa5DLkk+wy8UFe0ONMSqPeyfb2j5aIdpUMRHIsUCvG4V
JBkrj+U0pMUOuEZYUQVYGtxIfyDEikhHUDE53QilPxL/KTSZnYf9hEg6QAC+4Eri
SlLrXhBD1OL8EDZz2cmQaRmAa1Pkc/DJLLSLQp5U0iBmHr0XZeXagekU8bgoPabR
o/t12fWvPVsDKTom6zBQ7CwOXTmFtbfig6pFD4BSx6ROFKV7kptIo0UK5xbeBWap
klcxypzgVql1cTx2V/kLctZaIikH+2l4a0P06eQtMWGWwSp7RU2INPBZMf/yTKl6
JGXPb92tIH1Hz8uaJX6uRMMqCV2g9pEGHPxL21Fx79BpD+jQY17iIWsLi3ZcD4tq
6Q57gYSr936IBokhy9bndqDCXHxxAI7MCkJTZpEBeFGVhFv9WxXboudKT5BmkNAL
qbIN5KfCyjnVh2FR5CDRduLXHoI7xlt7pC/iQfiraynvXkVAgzhXfAYB5M9K3fZI
audvPlMeiVdd9DEAYYKcMxN06YWf8UdPrBJNgrWEhuqf15p6EoYPae1NK3ujcMDb
3qnX3qhEs/urtCpCztGWSWq7A/jzk59iYuYl9L5jlC4f+aDWDZtDXLMFqs4RhVYw
egs1DIQ3dJulyYcB0h1juZV0hR4feHKdaRi9xENgcZqMOw/Bua95HmtpmUCz+mJp
XWlAlhsF5rKYz4URJAVsnFnO+khdyuRgbrHVGTbl+iBA84/HXO30K9rm9nl1FKbz
y5VhhjNDPbRH5u2LgtLfg4qKtfR9rmBRrfu9GcvdS6EWaiMsQZzwoHgS3xgDx6HE
ljeRNDFc35rDJjt63oo/T1/pDMCttl6Kj7R6o8Sw4x/bbOhPDv4lN+NIwvvN6JWN
2XJ/xh3WrzpzZ1aNzIB+yYaN+UIHEmgVoAdpQNXmmyDq8M+egXbyHOHsaBi0BEx9
HbMJpQmgUaxIvXl3J9qf01wdCzA80ZRlMtHcY9dCjRdlW16kp/wUuAB8xyN9IvAE
wIUWOL/yraVKppA2uTTNJ/x92uQt75HqvOLUEPRrNZeCFNgM2UwVEMjzp1FHt9Yu
S9C/p536MLOMmMRKmDnCp0bMdledWWvDme3h6MQtdJlj5sjdvRMGvKd3UfRqfvdR
/oXrFFschmrEvdPoDH0vY9kKwFu3unfmStkNWKoqBB2no5IRsBba0mRnSoWFZPWk
/55/M3UJM5DwYx/bp3PlsAHnBikCW/CunL/NcyyOY8eN+jeaaNUhpUWA/d6Lj9X4
9BNHX8vk0adATRQ9W624tnjDHEaBB8rMaBZasd1eD4kcJ/JS7n+fn+yfn1EAkCxI
YpcyG272VUKXoE+ftXq2ccaiD943FKzpGvt5PN2TlkeEoTbd1zs30FgFc3tiJ4WS
c51meJPeAQR7aIZPuqB2r7Ok5dHORsJ1wuPiQZJ0Q4Sd8+puZkDO2DKTPtIVhAnv
Fwn6lmXYe5WYEpC+Bf+ibUMA6QrjZz+VVH6mPMsUa+xs6E3zAG0YVDw6x5TyLxcF
2QNaERoHlP4/s+/NT4OklKDgI4IDl/qIoexfoAopqZ14d82lH4VAeRzBO6NXW49B
Z8pgtcCrySsEvpzAip0J1wtbYKYdqcS6AkuDitzTwFgGnm37z7idXLadUZ0WDMQ4
qKzg1QnvwgFI0RqWnkrWz7p+vPjb6vMQF0BRP0Qq3phs+iWEI134OwXb6aQcXiMf
dUHXb2QoNCZ6pkf45yiJ1K9OPYQO+2mWJQqQh5LNzeEQfDyZ+sAxNicLF0dMhaMs
+weXVcFqyqAqvcQEzDtdIKzIznuLyduR5lXJxq1jHM1M7tX1YwSV7g+CkikJqTVi
ehDBMp/b8qigvLfT9e+fGwmFZN7nWBaXO7RGFOhumCZTWDHPiX5k1oNCcMMJ24VH
Dn1hDW4esqlBjj5IvXIFcKHcX/9TsFjb36tKiSczUxRRVO20MSj7/Vflot+TF744
Jm26N9d7Pll5BQjvXtIlSoAFN3nt9w1XAorJtob1r14QPUT4sPnfTH6RluQg8psM
r3Ykkm7z+zSJvEN7fwB99D8MvEsynCK1jNsiUHzkAqGXeXbn6Y5hELK05q7Kif7N
xiieHWbz+Yg84WCf4B3AytI31WnwZ/fFuaydd4iiHtkwtCLT3yTh6LX9Th1p7Xsb
gGlypmqqCPk9qE3D1cRszodJ61XAKKdbIR98Q9Ja2B/Mm3wgAR9zIGo4jRrPGL1N
g44lkI06gKcAfXekt9nWJkOSRoM15I33LyayXSkzhOlyFq5XBU6r79Ou8nXUMJGA
ie9WsuvEARNNy3FuDpBIq12vtERhYUo3HSCynAaoRcWKU1aGFYAckMC8zqr9pjsp
FgzrgeeJoE9gama1a30bK2tdyWJlU/QoN4prAEue7nbuZJmShZqt8n8ba2/nhrnB
Nq/1sXft+QstECpT85KMeK5Bq4bHSSK5OKXJ9DCAUJHb9MRgLW5Xhp9hf7x1RLFi
JrKVNL3RoltCedLNWsVVqyBT1Y6sGT8QWufb3yy9Gk0zJzNydlXTxnM+PRD1qhz3
ZuN/SGXdAzZJ5+mF/XjiilBSEHTqUA4KYb0yv8v5xztHkUtvs9A03LnSjKztGkEi
WhFp8Ff7b/g1j1ECfTP+y8k0+/qkN+Jtqp1eF1p+vPeaRgRPGmxRKRvRXPr+KDTu
y/1qh+WmO+5o1P8qLq5Z9Zv5pb/vEkbGjBDDRt3qsXARsaFKvo/WpUq9IWrdnFUX
4AYjcQ11CrcfFC2WtzWR3liyOowIeggUSF7qTC5uNjYuf94Zei1qaLje1Vfk/ozm
tpKqKrjVM8Hwhd79EOITzCyoRx+Tpoyg8cns9ss1+w1cwAlJaH5QxwN+RxX4dhrm
6KeitDrczCIgvnqtniBxTrvZCKmMBGGsY3vhwtaOMKfWKW/S5Pxtj8aTJaKUZ6Mi
fYTjI4m7yMBZe2XkSHC5DmgSAphFyRL6i3xElqu9LuAMcOkvoKyG7O9zo42bapfL
DlR6vgDMEvF2g0K1wOU6gU9ZUIdKDg+E5z3Xi7fNf4FAZTCBebfndEsW7n0GJ8R2
C6mMqfnHv3QSU3TgmRq5Ha6oxzYngz0Jeq6TVEgcEbv2dA00kPZTBHMptdXnENAB
6io/nOygVPHVdhIk6htr+L13vnVguKmvnewzNjx9KlSzPyyTa5JjUba+D4UqVeC3
qdjAdKN86ucEvC3A/7lRW1onWFiSnwmeh/3CazBr1Oe8CISYnUhEOh0IMCaEAEQ+
5jYFysuh7yG1II5TaoaAM76gVg38ofJ6uJQcskUGTq2ghvKd3ObH9a3CpAtkwA9d
FVLvW3LNwU3StL9q+M5+F0karXps6T4w/o3U/Dnd7HbXRiV+fSJIp3R8P9Qef3af
r95ItMZymNMQb7p+Ilhw7E29T24FkxLlpEc5KhJICUdozfOAk1vtFFJqcGdpgeoD
489S1ryL/ulAJuhfWa1ytCGY+ECSJMfh0R4VuRSRLyzmPMC1g53lKy1COwALQaex
VuPhnkYqqmW9QQUXNFJHvdPxFVTNmqeC9m7DVyUdmU6cMvjvwpHDbLVbY3YerGLC
90wr0di5MIafUvZioa2vOjSWTSy00lkqBU9Y5vkpDY7qn358fwt6OMz+cTKZDttQ
53m05ffruswMcWPGOqvTEw39qpJwhDZr10+1j/WaO0nytbq+6rBArbPu9FFq8bel
EZRkg42TpdRq4Doh4BkeZLW1g3IylUpDasOI0ClCu+VVYMzxOdlE3LVpN4AMk2Mh
ALDwrbFhqVUb4+ikDxsFh/tMCFa+I/tkn7NODr818Vi8541CPUIgfobmVSpqLsrl
iCApmsS5DQ4VLBLH3vXbIOW6U/toC2KoBRltMj9ZSh/JWZEfdTje4vq8gcyiKobC
xH4eOQ6j5LuN70V/ytZit4XJqATGNk50B9HN+cQd0qG9N+1NtBuntud4FKFX4Al9
vS06oEzHvDdbmUa4VWd3WvbJ4VjFdM3j9HPj4FEJuqaZRti8jbYg+I/ETG6iJYG8
FoBo3CTQlAemdjGlcIv6sMlE+aLYi+gQp4B9/sYOZwMT1wwyeGeBV90GjUO+I4JY
RZmuqfRgPwFI58/iVPIBjT092nM9Z8uDxufhIi2XO3Xev5OTLPeQmmwfLOLq5t2t
TJCq/rmK4zQzKvAQI1GRrQkcc1fBtq/3ueX82MrQg/phJw2gvgUwVhUP8rI/2h0T
SxEy4hbKL1LdechNcpCv1Ehrh0mXbh0XFXJzbn7ek7AsqU9hcsOG6gBAG6Yh6uDd
ZchQZ2inCzIrhfG5aWJhdMXXQ7/LmTwG+JUFNHMdvhSMFNY176fZWSKLdY2Zv0f+
FkJXmkXyOUbRZF9Edd7AXFA4MgKVyu0mzUHhyUrtga4ToMRqlltHIhWGX6WkxBkF
9sSdVhbkrfapvC66MiXEXAEFpgRhUnQF9ulQnCAKhBkB1g+Mj8UjgKdw3Kd6YuY+
ehxB7soTZhoOzMlRUvoieeTuiS+qvzNpTHQj2ABH6EoOvoKVoPoS6wPzzYzZhjlv
3UKBsyWHZAmh6T/8t0r6JEKBveQDIuRGHhVskE3UXzOlvHMtSlz6pX7QaORxekSr
hQs1oB7F852XdpTx1CBA1q3PxP4gOh8Foq+1dImZqkiP1Widw4ytyHwRGTFTf99/
jF5GRVE529zkfJJTFkLXnz/cK5d+cDIEKZDAYCXwJXFehOcSSpW5O0QPUm//JFPj
AhMGQlNE4zX93puyJEsRoURWi0aE9RK0hkBzo2vzAvaizitF6PC+F6d45kWfMU3R
JMG1kkg/C2OgcOuglsF+Ax0Y/m0zzN1dHN0M1nkhGyyYE31jBR7k8DysKQ0yCaZU
1z5uUzOvtWfmsSDP+t9SsspKftnjBMDvKOOu1Y9l+h0Iz2kQ9Rm+ROkjMUxKJFFY
KVQ+1lksmEighFa9Zo4SPdmdB/v4wYGpNktCTvillwyRzkCtYlNVXkzlu7XHiHlT
C62gYR4R24sl645nkBY5cCvCA2wwCc5IYFHiE2SG6vxBqYQqQhKs3C/9mj6QEadJ
b01ylQk+7Bc9jOQfvfaiDLdiqk4XvDRA/B3frZ4x1KmPuN12QLWvYEwQRhkJ0Uva
Dk7IZ73VaIT8OmmSElbg3j7yfRwiDL1A0p3ITYWEtiixmZMO9b8UYzkVG+JZfQb0
xFhDxkby9kcTRIZL85bwBdii5pqQMGxzn6K4QQAzlyZYEb0kyF9PXaHZW4cJggen
/xudOMzNVYzt8nq47YV77PdzyxukJSS+yaG7WHf8mvU+PftFiC98GNULAx79Fyvg
EE78ADsyo9JN/Uq79n08u8GcQ7FZgjv2bAjOf7VOp8Rixc/7TiA8H4JIUJJukmPT
8n+ETif5Dwey82WAMPDuzFkHpHqLBxLpotQNlRURAFQzZYY03SixaOJh21rv08NA
TO9s0YS2fTSG5ImDajNENraig3oXLcfS3OV3m88N+ivAA9TbK+6esUtq/QjmX7FS
MA3ebwRmC6L74IYB8EnSu7Bp/cY/FghwjdFGxLlIA8bOpypkjaTYhnfATmfeNYJI
8mr8HqJwyM87KIePECg1GggTg8xAcUHQ2rLTF6SNg4d7z0MCluazCBAEh2DROg5C
DNZXNFfjifUp++HSz6GqhLUonExHtIfM2GxUJO2pMaZDbHtAuiFhPd6I7tvgNnep
f1QxKXUU93w1njhbgucV2+UH/0C0stjIuyLEvgAke4W++LmGFJKOydpmpK0+INip
wIuE9C4iQSy7qzUGuSchPWAhHtcNXNYpXVKWkotl3zbAvtsde6s/OSYsFdfHkeM1
pb5ozuUuejymhgB8L3BfWbKeHdVPhASWnSjZFE4qFZjaPJU3mz0qIrsoT6vrdrnn
+CnPsB5RdZmKyPo9Iu+DFlARXUi9588VQQXM8CjnhZGjPnxM3kCyy1tz8ZgCyEXD
UEVcuHNj5rHNGjiKuSm1x+k/a4072NhZC7uVvVDpVGEeb/SYdHw676mFiNGOqDAS
QDq4knmil8nzKkPV3c/8ILO2OPRmsqB8LtAKC9X95mFx6PP0woDfIydtgqz0iJHT
oXHEXqHjoveYehsXztCdN8XxDI7Xci7GI37xPpJr7Z/FrdOOPOqZEQRna/vQCbTD
68ohvnqThaLVmAwUQb8dzGHWVJ1sRqr5BBXfSSWFBfkY7wHKlfYzwo4+J1eOwgWU
i/rmnDwHjXro/veTaTAT+lHK980uZTABFf4baYMAarEU6EEOb0x1YeZk5IHXllj6
mKTRB9B82/YgV2rYALQp0DzA5KpWc434IwOaSYr8FQ8o64NCZ0DzA3kKb95MUEdJ
grFw9Mo+Jlu4rlrPWigBHF+dC/1lZKt9vwAI8b4SdSokEJya6IKp174/7j+LyQqj
CaGJed0Ejs9Ungq6vB5qS6Xu+CJj1czQDPpHNO+wcPyCVhNq7PVsN21nAU8w1bao
iL5Uq1YL69nGGkrGsTjmLUU8H794Ofo1zJ86c3V5LDosHrIeWAXlyn9uBMJI8Gpc
aey8NzY5KIgIsLdj/Xz27dqe8JtTpY7ACqPjI1D9gqIft0T9Wh4fm173xsQf/QYC
K/opX8Rre7RJojXTsFFZeRyEiRmTSI3v7DFbCAEgJAMNRpoaOXL/s6JeUCkuyLHk
pqcDaFedvgGtstFrGR3r2O7QL885aDpeV3JtTfuELe+qAu+QnbUQM4UVSXNdON2O
EH8rwsWdWYLIoDYIsP+p1vUMEeX27Jb8tWb+qh3740btd4Uiuqp+4TmT7CKwdUS5
eagKv3Pds+a+/h+1mwNl6U9qStGusY/AYR4C6nqE8XcJfylkC2iHF/a4YrVkYKYl
PovTxbJZeL6hVtHaDLprUvGQtgF+Z4IgKLeHCP64Z3noF96EuY+1tj2nQtsB4fU0
xTuHxNk+R6yCaZIoXfhr6uC7psyEKxFq6esW2y8T8clkm55ocAbNkWXb1u4jajVV
DfaqJ7zBrCYoZa6AzpB1GkBkAnKFdosQuroGV39am5pm4qyI/QFkbmV4CtfVHqYs
yNIegFiqG7+FrTSGk2MHymZDhsAgtcr2Ns038JpHAIK7Ib2SOK1Evr70M6xqYmhv
ixsni002v2nLBvksF8v5Xi2hgzWpaslfduixes6hVZMr8xU9ED50RVI0/kbnPHKX
qIdR8+SpdDWDvgutr5BRM1kcxiiH0evvDD0NlESuWo6RxZVjor+ItbZwsMF+7yNC
/bq1G0hR+Cdh9V1AWMZHsRv6pnA5UNCSwmuIrbpirzPiSVg/K1D44oPi3/p1ues9
wi+A7LrjRrIRhrdWdvhP/ySb05n4lSncQtVnsMZ9sUOsocvG30AodVwkXf2/C5Q+
PHhXMQ+V/+zSx0b3j2mD53qdek3szM8lgO2s7aM0ffUsO+SSysuKXxd9m+dolDKq
fI2DC9bDrtd0CAiFlv5coy6RrUxBAeUib6APTC/9rcZ/PDhptx4dQDySfsDzlDcv
kVRn1zs70amrJ55TmnnLoOGg/SbiRozQLYgFiiR/VH5dXEtxXNQh5Ky9lkOyyV+O
shGCfZiZtsfdyKpRD6TnIWpjkfMtLNp6kmvqog+5TjtjGgr+SatVwFn2xQEkhjHw
bg8mgsHogcdnkA9yKMZcNs23XBJIFqyHc3VhQc69WXIAErhIK1oFWQdUUFctLeMs
bAeCF+lyy6x15Bd3Ctb/xEW2ZXOFiUd4+ghl2KHwSr7tfdS0jChX/bxVwxBiRV4S
sGw1kPRT+nixOYx+aVGj3zG/05OVKpnd+pkhTt+21tg/EsYDreLemhOqUACtZxNz
0IAQFZ23AFTNksGD8uo31r/ZXWyMQGSsr36Idvkzo4z4IYJ9NLHFeLGSwGp4cgnr
rDMyczLsRSthPCJxUzCFTvw+qmuuzpZsMtBLwJxpK9WBlcaSdgsy15eSn2tQ6hh7
i/aKJzk4SdEgL0JR/mZ4E97pXlz4G5mFNwnPmE24vOkNfgRCVXPutLsxIx3atvgp
glJkbR3OP+DUkEFv25Pq5Ew20SOR8m4zzzMW0HUXA2q2oAcEN3cdhWX+N0E0FnUW
vCqDM003G+PMDbIZy4X2bfKmncZmz30+i0iQUrcE5xCFGaeWoPKl4NqHPTp61fAO
361blP8akmtYEvDZ9W9NY1yntndCJXSk6GUe+nTlcFWwCINVdNQw9/+7wP3sSIu5
/5AJfQbjw8XxiPWT+3wrmIfVplL1vdEUMD0FLQhVpVJTt4+LHzV/nOoLlzbuvsxm
bTWcJIF2L56aSGmtX03QA8MN+tIIyB+zSlzpjlMJ6hNii6waNKp1X4+B1WcgoI4C
YemH4rOdfiflLj18dcQSkTCbCT5t1DU/UR0IMAYWpa6wp1g35xOeODFOyL2s8RrF
lGpfmBWlnAh8FLJuzIAnbpayReZqvH+ahWIClHkBqzQxtkpkA+XE5WCtLf1EsnkS
HtYXoSdsMdFdTl+382eY6MTb82262P24NBrKIk0mddBqX2HzGrGqJq/GS/wIxC9k
7azB7biJGb+6QhRD8zUj7UukGA6T1n7B1HSFu6FTU8j5s9yPHl5ZofjkTxVZCjZZ
qWoUdlEoKY7A2leFKxAd6QPt+JlZwyXtRxYFhH/FdScH3W66CbG3eD6urieWCbdz
pTgtT4m483NDX0v3ma9e6TalmHkbmmUKF/3rKNsB7FS+LCBYgHLhgvc5U9NnAnJr
qhKcntLQlRUGDh/PZuXW7zBfmgXvEaxoVg3CMT5sJyXLs/XmVxw1z2nmcvxqWJ/d
+zk8ffAqjyhy/T/joL5MA8EF3yo4uD7aln0ynHrOyP/NqHSBfbFWQCpO3PWt/EH2
dTrukVJg9elkgIHFkamqBW/jXXOF9PO9u4Jmsk5CfmIX5MOu5MYKbWfgaXqroYKZ
BrdHxVEnd5oEH9HeWESVqy6IpoIry+Opi1LTOVpdmocns+E0NTMCv2gOzeFDfGxV
g8T54S5EsyCLzhi2J6JmfWtxEaiLcLNCgyOV6kOrbOzeXlHfuf8ivgqucNDa/E9Z
ewPYo8UPoQEDLKaEUWsgNOv5QfUTMUyDCFJecRO0d8RgyX5Aeq8PWTXeWheBKXxv
gGiwltiwNx+jpr6qm5jJnbQDbDKJzGb4Y+s/kGX64sYEdrTQAOsCt6DJtwaUuepZ
KgTV1lscNvnCs3/q38+3kk8ueew1hN8HmbAB8nnwAaqD3TorQ+H3MbigeQ9dbMGy
BTo+Dz3lnAxiYecEPEP4NFfryqdB7HSquEo7KLGWhmbMEMwdIjM0LvtupFF9qbV0
/eJ0dnN17pJW9xf3aPx9L8cgqM/jqDD/i6TFlVymVz12qHuwU7GvUoJIZ7KyAFQd
qM6hIJ742Y2bru4npIVofzY/SERWJl9dDCKK660iOzJY3JgUvP7kfKZHIDu0XRYL
tgCh4gV+P55sKSHxggBUTpzanEwt2k7CoN/GxR3tL696cXEzBeEwTMmXWfjHw/Fg
hdRDHDyO3NAZ8SNCKo5i++JMbed9uYDq0yRvaJG1y3Wr03hjGmDt4cR6Scw9nLux
lV9SyB+q4yCCwHZ19OzA03q1vGUsal3E+WaQI0Jy+aUj+iShAfejDGgG79R5F08b
6wYjuMm4hInJtI/f0tzzT02bvYaqaPPhuuuF6S9kjVye1MX8/JZz+ZFU0pjBUpHT
uem0Urj+HmzmYLPnLxGSitqbjQPb9NKoPVeDMcsKA6BX2/AZhIE4Xv82EnYNiLuN
Vm1S3FDqZ3zAerk3jc+8nnbKULiJbIAyIpnmXJBVniAlWKRkMDZaJFWlhcdRvCtu
3bYxerYxE7hdlTRRmE8gTGWF+o1uYj5Z2s/DA0IRXrapaQ6ei59MDxPlOpuQFM0O
J+F9647W0JC4Juou0Qyo5EAhpsAGPQ+A+DyaVnBZb/hA4oMJNPXrJbUNU53yA7cz
+q2XCdPxrl2Ym5k/dqFV+D4mGveclO3kV5iSYyVky11dpTE+2cnrP4fkwZkfomRg
Zw42mfjA+mdm9ndAwvIdGBAOuOMa76fW1e8cYQlUbocIImYK8BrUWYjavr5qiK4O
W2YX+eOLoy0ATW7uTdEx2SVudLANZV833/+pes281Q8oYbT1GmUl5gnKJL4xxr+x
5Hl1O6uuC2nkLjXi9sHATYbtELWdFG2Emaikj49mW0LXafHvHGmtIjiTluNLqmkg
4hirOYeFvP5iaKNd4rG3Dq99DBVjsLH4mFqGFQgynpSo+WsPUiiPAGH+PLUN2gmB
2aaDFC6YN8r82/jZ8bx45kYTHuDGz6+1jDLXnebHs7lAHRYzUDsThoWbmYNOzRIt
zv3JlNOO6fWZ8qidfM8o8KIvNQpi9GWmzCJqEe9pFMNEw8R2sv7pyxkgE80rdm18
c3xJBEcHh+uX+/It5Zg32EGzDkHzDX89IBu5qMWUAR6HF9M/7CP6A80Q6TUbG6tv
7BdpQ3cMGRFpqDjIUXshePvr6sIsU0NB4VZkLsODKrrkYPo8Q7ad2J+CLGqqCZQp
zb2FRGcDmdocYLUdBGBNt83D2mpuneagTjiz22VrEtThT4IBK/pIjU1+Phf2zbz0
/1HCaKX3HbzEtgQYjwAZVgwFfrqkGjkCjusJx5w84TKXEdwqTUfRAlEuIKc8DP2F
uyALREQrfYWUNhRG4CjwkhPi8G+CLZxb+W/CTClUr/gxqSIo5Kho+yESnsuRURdD
r6DXq0xFC9LEXKcVm4qmImBwr6odouGfDbEelbV1hBhukujRn2AXzeIIMKN9fhVO
PCoeOFywa7rimZmDfEfpSXK59teUJo7c1cagagDa3qHwVjCLBFmV7rYbz0MRtHVG
GrwR6z8QlMmjmxOGj3b4/ZHGnKp61ISyg8wKBih6n1Ke3oM+MCxVjtOh1VPK1jCu
5+lAKOSHkrLppp4p3fPmZA2bSIC9Du+HMtC18X2Wdt0qc/owD7gdEp8Te66saFv8
6VvJGs2ESPNTWT6tasbJcd4758/CJ6oVKZy/tEnOC40orheEMZ/QUoXsYNz866QI
7MgvedeWCLnJObJ9hXuvDKSYdkR4FSI2xmPXRXDKyd5Dc6X/CAWvqudWeeumeD9y
lglFeJrM1Q8+FTiBu4zVuQfLu3Dzq5aNg/qYKUJB+1SsMp7ABqtFYDRGkrh78RK2
n9bhCdOZT6E0ltulJn80KyXjU8mqkKaEwpR+Y2+O0ARGJ+pQks3uUd2oe4/TbWES
8yzum8RkownLgYvkcTLWWw/sliIDIX056aHe2ujLKF5Dw2i2U+ICA4Hgl3SFf3vH
E1Ihm56733McnTm1PlH3drydcwL9eAuqFEpi1ncecrPuzmtZhrB4/x6c2ByBXHV1
bIYx+YkzfJXY+YppwhH7YdVE94Bq3CQUnmUvY4Vnh32feQReyjtEUEq91JUbUm/H
5H7N10tWr+aNdhm80AswlfbOXJoxhn2qE8TuhYj2DTfLo6YkNTH7h+IcaMQq+pNV
BKGAHZxAhrtWEgdfQNuAK0Vv6rFu9CAJKIc8A1XyqMeBYz9El274jpIk4PtLJow5
zt+CFi+W+rWgWKLZ8ti4pSm4JHpirAoKAWaDcvoN754JpLwfxN0UbgOZwa0HHu1M
nZ76H7TTbx7KldP9CJa1ZTWPFjokTyqEjssrUOMvHaMNP5EfT2bXSQRgP29KNuvr
HokAfMFaARCHippsEQ6aJ5s8glEtLkJqKjOAiklXZ+oQHm8EvTzn2pcIEmqk+hMU
17dqDPd54zUHNoE8dLFdCRIb/xV80/gNsb92V10C0KNLM3HO6EesTj8hVw1/KrpV
3fENV7fKh/J0xciWIQmEhMSev9l24oZaLGXgyOzs4Cr8zNqICqSdwH9OsmpZJvfT
A2Gmu92puJg4SpHJeO6IWIarJ5yY+Sl4bdMtokQWyItE8yuTb6PqYEgOJ8PaqJcI
2N0/d2scz+iFkStZgjNFhGAR4JqEG5LBnkYbRHg6W76PZEzBwXe+3cb69FJaWHIE
/pg7Pl0GVIwvpPxFPB5B71qvo8fDnbjlW20XsDXU/XZApodoDl9uvv8QAVfyxmUB
F7jyKYfsj8ZXkXod8/kUPvIiH+Kr0znqLBsJnFZp/x+hFpDVaCgCOeAutS8wlj2L
nfnYFvgrujmWKYGJ3U3TP8UZO2uOU198Mlh91qmpIWLnskah9skq4m97JixIe2TV
NylhMC8tE1/L+DV0Js+/oxd+RVlLuoHZLnUn0pxCJp4ZGA3gNqLu+1rv7I3alwqq
iivVSuyBz65uHtTlR8xAw/Buhca+/pJmxZCkbjyFojea34jM1C+8ImhfO7WK0W1b
CyIQoQO/a20uqiBHKS5FVSgd/LO72qmdaOSt+WP++rnHyyMEvLp7/JbFFMG7oKia
HpAjltHRNIbEH4n0nE07kUNaR1sFEFRfWWUvqMw/m/3VJ9WI35qJAJ7QG1vuFIXe
bg2t9nB8kAUzFYbick3RPBEdNatmLPtQVc5b6IEVyIgLxXS2iK0aUh63Ep/uXaw5
VGWmh7SR/22Y6g7RczCVpTKMmuoJDXvDDaJhjhIRhrC0XEJUgllT3r65PJWwj/v4
9FeC8mU2wzVVfX2avbEXNgaIT6CLrgaSuCqXHCHXAhuL2v5lQ9ML5BmLtledFpHs
FPmZ+2GSHtTbcdu/ep55/CJKMsKVqer3mues3eq4n1Klu5qi7GxumcYP6pBG+VLK
owZaP5Zv5eLJnsB7ZFE9aVXFRXRoQCt/aj/v/nF7KGvEmxCNWPi1p/vLY4zcQ3HR
6sJEUiFKHSWRaZwznrNxBsUWEr5B9Uq3A2tHVu51YiUwgDOSeezas2Y8CNPat/Si
Vd747UGAqQmvl+hZDKNWvd0zfk5bg0+3EFsD0jPvcWVc7y7a0LUbOu7D41DbcU1m
ayaIbx+jne0eLgAIC7W+/itCH5FbRC+GdNb50zi9G2UCEf2Ju9KqBN/y0m/8lOK6
jhmynOpNMNYBIM29vXkDGfcp65cKayIEu8Ogx0c3huk/MWKVrNyH65rYF2sEIeYz
lGlR4jT4ncQsNdPKtECgR5DFloFn/MtMwwW7PnSHETnnlF8MC9Hihrvsmm/2AK+S
9h72knxw+8Pn5RcqObQrIPpKhPhXwTEqg+KdTfcD6S/bFX8iKC/bihsaxQtaswnC
8gYf7xbbHO0jdo91W/a21lwC/1SPVysMFt8/VG2Ie7PtJvzeEYsPNp4DmV9UEypl
kAKxx2ANJHgcT7/NeheAq8nLRx5pM5uf0B2X1FuEwdIJnHN2/wwjzsnFY+TbD3+l
1LDiRKlf/CPORqVn8INKyEbQ3yIj/w/hbR/TyYHgrY29ZDkCicpzfYjRoGyZkc8Z
ABHsM2YqtLDLIIBn3Jz+tmUTmzfegIgAxjzE3tY1mAaFn44WRXVbb23x0exL+G6P
pVUt6tQ8GeXzqL/MEkntTZoTsqnj9/303UKqim3wZ5Pgh0U12eX3ieiCECdX3Peb
xOQwG6kTd+Ss09vJz325bhZAD+W/Stx4xptLAHoXxwEOw34LX6XKZuwT/3TM7iuS
pMtFXDdTFgWqyYXCNVkwLohw9LJhO4OhCo/0ICkZpgbUw0UhnxcTtcnAgAU02wVp
o0l6zzpogK2xZVCtUysq6urMG2UZOL0CGmY+/X3TASFQnzHjNh5Eu4ukZE8xQhf7
Msxyyj7aeZeuhAz0eKbcRp1R6tOsDRH9lgaVtj7m/jo57Q8MgpwHunU3NWsdVpzs
2xa5HFh+YU8++5BKRig9lp+k3dfPjpX6isefXaQ3ETda2Z3m+DlkZ1C/yhRVbcFA
126X0fX849uuvq7xXuiwILD7vdFbmcA25RPe9oADZ/3Q80AYONMaADUWuAahr8QP
uQWND7nfuvPBa7tVjgCRivSqPwGzpSvGJgdSt4dmOF1PrKbJJ/xlICB3d3aBd1rZ
C+r0w6HhUR3Dlwou3A2v75CcMP1X/DVTO8Ue7wtboZzalKudS9hPm7Zip7q4WEQo
s/u2cdH1eF/slbFXWQQbLU9+v9Gj/9Iwy3Nr+CUoeoNs1EhSwzg3gSJlpbgw1/1b
qEYnh6OfLyaWIKGWyGhpYHiA4/Vq8V3tqg4RivVBjJGsV0uEEL9no1EHLLXBXtmW
+Cx0PIM/tr41RWLOyYFsvazNxOR+MP4Yt1+9oPRVvwysTIR9etGl0HszvqQiV82e
stix0/1oO9dsXVJemsEFycNwPZ0qEi7BUUdeMfY2hxd2xjYKxW2LQtfldMMkmdzp
bpZxieYAv+O45kTxWZXDr19wwXYx5EnACxRhTeL3+H7ld5ZR+HaQY7yJIQDQa5Qv
UuNZ6s2gckBW9qhogDEb42TmRKo2OAVCZx2xR4k3QsOZfXfEySMJ+avj2nn/joLB
iW3jz2rgumwTftKLk6oL8L3DU5sCuor8sFLNan9rxB8wK2/dE4FyGqInCuSMbtmI
DOqt/ZEAyquFpuvr1zjORP59PX2O63fgW751F2fecKQzccbDbWfJPqlG7YUQTWLg
1+d8DYoxNLsn1fCykgbx+YFyE5d5D9VBJfXfR8Lncw/dM5kOS1ngrC/13qg3g5LP
0x/6yOJ/PVWX+asb3Z02nNE/L7ua7l7Vn0/uAnERwS4k1GwoPRlL4hfp6dOo68bT
QuCKhemWrE1COn1pmN5eQqMnCcC6+Fe5bdroirBzD3dTZyQ+0ZKOd68MsbfM0WTL
Ov6XUikRzjjpZs2G9ekEi+aUugcojR037bFxq2K6TVK4kMxmwbAPNpxSqBQ9z8Eo
3QtvD1HlkW9YTj5o6xbDSY8GxGHym7qMaGlPeTuorkew3BlSf6j+CnFiVdIUEMCK
0pPI8Tdwh3iO0plE65nKVbFPNy0sDJ1uyc5Lqj2L20uuKOXNNHm7ffgoQjeAvls1
i7M8ZbAkEzprrmgbhx6PxnURVDHFlLdEKJU+g1gKJN3lBD21GA8Vga1Sx9zB0oTQ
cp8pvu0Sd9TOHXXtcli7JyQmA9JOzezQJH+RUqqLAp0UDX+qUZ4Fg+lCzhTB9rNa
RyZ569NdCl0QCOMoLEf9R5JODiegd25I2HDUpLNtXlez9KaIlVYa7cNtuRt9ehzg
s6WmLdUB/oXTVfyKPAS6uH4ACo9gq70IVcaEFZDtjXqlf7IRMlQF47IZg8JeHHWV
QD9Zd4tJq95RPxQKs48z7Mx/Y4g4eST5St8LBXh674ZTOzelbQjZSG61K/U8uyXG
n0ctpKU1dne9Oglzso9jq0jtOwpARvQptZBQ/jZMFCgV4DSZT04lQBI0kUeT3KOH
FRbO47F9U7eexHd7XMPoMJWtEbmVpONIpWgmC0d6fcRXnK9zAg8MeEtxSC+0Vx7l
zj2dSP4GDXDLXOcxpcWBpBKQgW9xojs/ucWN1UQfC8M6T0Ya86X/j0NK1MY0VW5U
06IMqTqgPJY/tlXFb+S3axcloHQ7+rs6IrKNZFowKZs3tN6MeLG+vUm2M77hLqeu
bbcl1eigZK9M0xLXZy9wyHKZtr0uKcY2pMIk8jaQjlhIlcWMOgbuFGtpddauSL4e
HGfnR2bs+JKbCxfH1BoGb5HyWbjZRSe7iOg3sLPEQJaiQ78qm6XxcoeADhTyJ5oJ
GmuJCWX17gKg9X/kq5TQBEn7sVwDJOUMzRI8QCpe2Fx+58MuoyAXVIG+g9/HyQOR
9HYDxxqf4vpqL4NpIxB0mo9wbvb50xTX8BJqA6LCCcc=
`protect END_PROTECTED
