`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
O34VciC96xgpIoDWkINKVQGzzIVwlrcpWfynBnR7ZYRImo7gb8gfRGTBpFeZa9bN
yHiFqbR4kg7cJw68+kkmpfZuPWVHnRgJ2rAiLEC9gAdfJ61gmZUBBmTOASDgi6rK
fX8rC9xEHvZbpzWzDUUNlC/i00Ne0OelvUboQfElLMvth6ITSeirZ2ibWJNLTy/9
+6X8QuvJ/4VwXCh9p3dlkYIDe82Ax+164P/26WvESU9YJL1o0Z0E5XNuvpxiuNNb
8gBUc3hhU9aXadBOUmHlHHcgIjZgtWzlfG5sqxJguqx+ekyMZkCn62EZAWnGnQOm
ZBaNAS0uavLaZL0ALsYILdlPrGEp9eralfayzdU++oI=
`protect END_PROTECTED
