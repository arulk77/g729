`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
sNuRlNg/I/MzpNsqliDkCNj1ui4oAU+b0kGs5jUhaEAeth7e98VYzm7BR53DDVCc
KILlZPev3db2fjBgsymLrOfx2h3+Cb7fKukv4QvDjf/fMyk5nYSFAZ0V8kme+tYF
rCamVecvEyTg8qbiw7T9578svDEfFyV7jkhgmY1B01luiZLsUb2FBEozhlzDnO6u
Pm32acHnQelciVBe4XQ19Fm0eafuGyLPakdaCBpg0JUH2Adyz1jWHShA98zdftPn
TOVOxWN7vpxBuLSWZgvfK9oCYezdrPxvlB3IvLxt7QGRl7JfCq+29FOnwIn0TSuI
hbX3wc5BGODwMj7WRo+adPvxJn738y+vlh9JwvfKuXNbUFlRNxuEpXzma5p9l2jN
sYif0j3PhJsMRgO5Klq67fEsyXP/ohOIBipqd4F1T0/OmgME5R4Riw48GOkBxCc0
UeQm4Whrg3nJQru20DbfyEbAAYownpBjgXJba36GPf5JNnTacd5Js2IEvgLzvtn2
N/CJcRoHthfLhMcnfVGnRQ6XUYwzqp1swmtKEHggrS6ZYEKYSwsHnxmeuxi9Buzf
JcxOwZYKzhKCUIswW1ch+Qks3ZpFLcNjujk4T8yG2a+HGFVdj54tLPUnazOtTCSw
tGefFwfgF1kJMOiZUOy2QI2vgbrpUtN1fHYghxp/QWAtrrgzD/1mKmnmv2g86sbB
vZS1ejqx/hkrshQw7bMWSES+lJ3ybgaZZOlRygxFKcylcQ4ONgtS7UeouC0my/la
8ANctp8Jy7Jwa9bKG4W8qjO7fKo3rPIQTL+7QWNojEvU2Ydlk8fy+fF9833x4GvN
fTlhC/D9YXn4wtF7nsqXjg/s9tS8077qHkjkYJ24KsPg2Z3hKIRw47wzoGVExfGt
DoeSKyzO4ZsjeOHKGzjHNcx26nJbpEXVFvdjTLFTdPo=
`protect END_PROTECTED
