`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40TOeyvIxRO8z3qNJNMFrdMNgmzDRY9QJJp6uEGiWB1l
2bSk5FWatM8pR39Q3u/ziHkZTY5U1OUXSqHcqtCNM6mH2YyZrQtCLUlDx+jCURQ2
XJXjDDCNwdno1qnUnXTA+1R85gl41Nkf9aj/5AJxbPB3Gvur74kd65lm5gct4dZM
nngAkyROJU/umtrGsesMfSXrHk8fzWZgHSBUgs5XuX+/O3OlgWz00MnjO3TBGrli
+aDrZfRbuiNe6Z9Ku6exYwS3zRsb4XqVoJx76UVqHYdizpPtgjbNmbh91/N9Ae/x
nQMVSPjzFRr9cbz0U1jyWK1kboOdu+/NYYE9GN9S/jye07qHNpGhTpQ2AsmiNHYe
S/+0wxYCxu0Nd8PnANf/r6vC3OachqE51wN0hfaWMOvAl951H9XaNv+JsCuDSPLh
zzTM8QqIrIgVsIywHYZPng==
`protect END_PROTECTED
