`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zeIYLc+jKW8jeppYyGT9pX7crnVnpj52ZLSf9d/2Kpb
Vljts8gsiJUdtBAgWF2TKXqAqezsp6XKXHAKMKP34nnwq3kSpjEQJCLrH8suY/uV
/BL+1hLK2RF0h+Zzm6gyAavLWuhnexUJT8girTI4UT1ngIrhE3gGXyJwPfU4G4Uf
ZemyYkiyOLDD9K522EwAUqlsJwbbV27uKtLl94jJd1cOvHBATGPWeKjS1sJo4aQN
EMxdOZklujHibb6Ijfv0qRRmzYqz6hHC2BRnstFj0VFDIze6yeg44XUZJYLBKAsD
WKI0lIIGv8T/x9Chs0m+S7DB1l+FbE+y/B99gh/9hA2QwexiIfJROTD+esjeohv8
D+WHNphTq8BU/NBvNQXHlQ==
`protect END_PROTECTED
