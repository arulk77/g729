`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNC+mBFVJB+2YdZJMVQmBngiORGcC4inNPTdAGq2848M
elpENz0dPJ4fAMKOxk1uKEdIFuanawDJa9tCdM8FWQd1HFob8p4zcSC+P1nDQYeF
tdEz1GaKyXvq2/O/fMWfBRV0h+67fXMbaEkNlshQBXBE5XLqXxceREPY4mN5wNiV
xXlOkoDBHAvicJuQymrcCV/Zk7Kg5eNxb/jm5fH/OetARzHtbGDgnqD1k4OJ8eYh
LmsRUbbwR+zAlZmUdjFjUL+B1Dcf6SjWkNzMOXgvIzAKWoSwqPDrOtBH/QQVhPHA
hdGqE2XrXZyWSU2g/KbbzA==
`protect END_PROTECTED
