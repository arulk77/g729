`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zdfXpevyjXEcE/6EphnivK8BXX20KN2bkElSyYUAodsiGI72V9i6I8gPmw9HFTN2
pIObDhaQoAPikVoo3oilh9B9xAE3EOzDkZNwQw1YR9SAvLUFB2SXihk2CQKM7TxM
yT2Zq4BiJDWc+LjeRv1IPXIK7E3UZJCApwuvNvADxbAHvPHXJ/7t00Y3xEZQK/TH
Z/TgVt29i7cT/BYKydj0k58gV1vsaVjBjk1u+u8CVF4=
`protect END_PROTECTED
