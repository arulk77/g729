`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHI0N0wiUGQ6gyUwbaOoi0jXv+k5AyDOloUli231Fics
GEbQJlb1Ec6h/xdLUtM7ZPUPc1KbwdL54sdwFKJ4iSNuxrnA3oW6y1knJDYDs+nL
suoQwLnSctAJfTCLRNpVcywBwhSlImeLYYjzKGwcLdfYARFgvVwtzMJmR442NCsA
pVKAmHWKznjlsJsLAmg8DFEIwgDFz5QHlNVD3ONdlgL5Br/fHi9aWPanP9DDtS36
FmxGJuYfnxV5xAJgdzyDi/lK2cxzkXqzn9ZAfM12rDis8qi6XeGHtWg2agarWroy
Rxz/L2+W4ifP+ix72IbHm7/u2hr1BQiQwi5p8Kqamrl1BvpsylmnDljyAWUhAHLt
mTG8rc7rtMOYxcW5hXxoYmtdAOPN7ky1IVwRA5bswcGGzkvVqeOeq7geJ6kzY8hx
xohLbJrBiF7YaZx6PGgh653wsbKBgbvQsQ25ad2sez5QjRtfVUw+AfGGiP0uWUYA
ZR0ka3wPGthNtIvx2R3p0eygttMn294QgkvDCFFoU2MoGVvnHTsiHPTqRDo+AbJn
Qt7nKHhsGqOxULxFtUyjwHnr1ol2QadBI5mYQXSVsySakMmnvX7X5mhOhr5izL/c
HfHdJ/jry3i6hLX36eWm3ep+b/Q+tyWXDFJY/l3I2l5Nsodm6sqb+5QSx3w0ErFp
ivlX0pgEQ7zt+WNmW9miZT1/f6NoZxk39k1X1Zm0joMvTzmIeIYdjSobNnT0F96p
DBepzSL80jkrFw2b7hN9T79Ic9U4wOnS1Qc1a2QqaQbD+Wls4XPx1GLqdznnmC/5
kPR3kpqsxcqBnOqsJ9RbZXWqKzAh2dH/Q2fkZZudGRIdBcQ5KQIJf3C6+cIb7sZZ
60qdGXcaw1wMVT80reMyExa8rtmgGVmWJNQZGX6YpKq+xTk+Gq8YzID+dfSWSY72
/ALO5eAPpteIYFXzE3qPUXtU3r5wbUdvHSl9LCnRajojOsQpThquNKBCAjTcPaPh
WHr8obtDTYD0IMQzgywBfMh/OeQM87dMKmWYRBl5aRVoq7I3uRlphm3heES/MK9A
OEFANe+oaawiH5oeIEULML7CUVfT9/h7JHSwHUjHXFydL+ul1OMY9tjK+EAX7Rzk
Sf1x+gXdgHFnAaKSBBMtSe/7/uzJlRZ00iwnrTsKHK4b5I2R4ecqjNh2M4NY1s7Q
J7rt5AOWvBXiMrbFJPMLpYpxYHtF9LwMl9J9PecVoqMQKy1qcCsFcN4PzEpSjO1z
V+rtLgAYk7fkrBwV0c7TK4IPxXZKgEsJ44AoDBC1SWjeQy+tcFP3doV2fIod3MNz
5YXlj4pFqEcH1+x3M0NhjvSZbrLSfD/QFm82LRofjFI1drGnW8P7yyZEcDH7xT1J
AQJU9TeIVw/r8wZBMLKzQMUW9+Jk7Vw0pK3hv5IkVWvyK6oVj2FcIn+MhO9qVy2h
km6KeyRoTiu6X4km/NRULOkqmI7dm3E8u+QXK3HfovGsI1NmkdbithdXkfRDoIjV
M7KPvlBa2Gu7lB5mDZgfBAKTFv7xIPdFHihlfQ+AAdO0bCqaoSjvEHKYFahSrQDC
BxhF+/sFj0FnXchINBAwODSfe0jgS1ezUovvft7C0wEVj1E2WTjHuO2ERMfeSgoN
X/zIL/yA09OMsUv0ZZhnqXHlhHN5572X+1Yd3w0RMmbjEvTqdhDjUAfPwftuvasW
wrgNmoaYFRnegaqSdcN4fGcChGOOFYQD7wPeq3fJXlCkBmkOHgcnMdG6ztt3Ag1B
5qDsXDYgdxax8NFSAqt2do8OmC1LoKDhYEeZkVj0uTWnEYZMq5KpldkOFruZiGOX
OFJS6HG5XYtg4sbXkFFdfOcNwqj0XrpNdYUar++sDh6xmkbW8sFwVejCFY35TY4k
ywyIMYu588r/2ql6sY0dtKMbh2ErTlV/gWI55xzvN1G/U7uvmtIS+MHShpn8/hXh
byQ4qDvjYRmNnJa04oyDkD74NSMy4vLR1dOr57+W0veoPlItTRdxA65sWMkNtiW9
EnucZO6FyXz4mdeo7QaIAPC1CkbHSa3Uz/Y2UT6pLe3T8YyzPay+LkMVBaMepM4X
KRpYFx0l0SYO28gkA68MgDguEfGgTR1TSjIRU9l5iDQnMtbVc7+FxwqpkvJ8L8FW
TXOLXvs92YuY8qDf5K9jQYv/iJXhrwDTV8TEoRLy8qHI8Xjzfo1/ayFgoQ1w6FYL
k6huh1+w2z0npmylc04o4QY64Dosjpnihkh4we4RVuh7kXyCsl/aOjtGwkcdhBrx
nXiktiracdi50INLbgJmyrnKE0ckoGcFPEYv1lshhYfY/N6GOoEemFQKBUYMh7hF
uN+ZpJ/vBasfifB3++xvb2lIDuKjIs85w7IRSj07RCv7ImuwKg0r1jPiFLCK3LoB
ejHelud1P7/Q4XC4CAlg0Yx6f5eT5bYm7wGqd/6ZeImReK1cJQaZHFJu8HKcD993
yQp3LeVjxvquZidqnxAkWMG/x41UzeZCQI8dUjPeiVewYkJof+N+y1RotYj9x9/r
DZfS7Tvfe0cF9yNHW8DdT1BtHx+X87lxb9jseyG3q1mmqBcCulbA39MHeGoKkhCP
3iy2fAZErM/kuH48tVK7AedeeV1ejVRSc5/HzxTjrJzn019//DUL8XfmhTN2vr5K
iSo+G1jaaswqfrZATQlWEJqD+Gau4KOXyAELVyfWwYPMxVyCsb6rtav1upa0bMUz
/BTfh1h2Ha21uMuyhhCWgQFQrZ5MNgqnm+Hb+yA+lgzklgh0nx9D0GrIR9vj7uDO
2XoNuvl2D2+OtREHvl0b4BpV9FRtrNB8FlOiQYRlQLA9NLUh7hAe5QBi8J58C4SI
T5et6P55+3+cPRFG0YWo6cxx44ZeV8DWdMOTunrSV0sPBI02uD64uhu5zcjD6EUj
9jdl5YaIhVSgJ1kOsk1v5+0C1MrTdky/YTg7VjFCegQ5utKNDxw4qQ4Ig7S0PyAT
bjnejt4aP1wUBbblYaiLGRN9+gncQNy0JykYIR4BkPHAtDcIR52TS6JmZ/6Gg+Q3
O70pQVzSvZfxHYobQXAXQGgginDbw+dAReG5OM0TTagftPXikPbJcbwW3XzpvCzR
UpkCcqPUTRuA12XsO9G9RZ+MMXYqmJZaMNVeW/pm0t342jE51n8wp01qOoHDDMQd
rIk1PoCDsM1sB1+VkEcCTfU7aloonyxS/CJy0mt3Li+dSJbzTFXZhiOAlWr1Pnzm
bxP3na6Rf9FzL4C0aATHuYlYqijxMgXnTeUsiZ5QJz53rU+0WBy3WSDD/teiNeZI
Gok0Ko/RlePoRiWqqFhcnpUnCRxz5eP/45MnaHhbejgSnRTzfUg8ooL0q1mSKKSo
DSmSZy+u104LpIQFVOYeEalrnaw+WB0URYFkgie9+eGXt25oNEzQsaiFq/6x2njb
rD2Rb9PeA1+A0rhfQxqL87GjBr/k49+EXJaxmt7PacFmHjYpJ1u1D9aVmvYse2Tk
GoVsIwKCMcxiCgY6fAKeT6LPkWOC2t/q/vw2A1nsn3yxrFQCiI03M6gurMLgZT2l
GaWSO64pf4c+xuHTsrspUf7WWtVSA2Kpub07AgZNIIygxIbxardegelwCXoKVKks
hiBBgFMCf+CDjty+5HwAi3mihYJrxcXOFVaG9TkDQrny+kNpBpfYmw9LrMaa3jyv
YqaYJl/3BTv6/xz3cdJbw9DwqJWA2/V5hRvM3vy8mgu4ePD2eUXcE/c3B9tOA3Jc
GKj/2J1YtHNt7GTpo8TbwxyO9NmiRQzAXSM6YdSitEVv4rUC0p10A1d74FWjUXxI
6jba53ea3gPxi+wSTUkGtY/5HoplbDzqOulNAjXQH0sC23zYqMeiD6arf0iSNvn7
ud2dzejRu8ANNosBX8vOgcDL0e/OStJdtkXEnkEMv/xgw67FvuXo1KsJvGx3MGR0
HSjUXDOvzPEEomgmsmNCfdM2k2mvuTljreGjq3RXfM+qq1loETay6gVNyC4cHWS2
XgRjOxdXDcwnqF0z7y2qsT7plQ362RzZHsTqwFSJ+qDf4CaEotT8JClwuI8IBgQR
sKG1xc6P7gj63kYB/C4xAPROmTwYYPmgWNAQzHCvk8xeM1fMsfMMea+MSgKC8/YG
K+ANVUviALhY7BNmNMJcyt2aSLUqaX9sdRp7jkablQKgvBwK6AodeO2NNOCJ7YdP
raGFAaC+7MhAm6IV1M27a6baUZFb1JXDLmGR8zfbnm2m1JTEZfMrrwMXvLC9KJ3E
1FJeBCz/nIWYXJT5IzbzcFaiN0vlSd+17hkD30V98S9GmL3q62JMm/ndw08Lk2Qv
UsE0Z0vMKN8ItiZca4IC4YnAYGGRrxsy+lDCitGDPIivGWusZB0XJxQqei8uhKM9
ZBc+4Qh1XQLEI+sKKW/B3fQWPMe0LKa200yJrZ2SgfZuUNTbCBMNYJdZBhToffhF
QhfmaLyZhXAe/Mzc8q18yKCnkv6EPaDd17hVRXJ1o3zyjrMJdyZobYMKAxuXodGK
7CxGzX7NFqjAGp5t1sx60v9RvLsB2AjMvZHYzbGy+DeYFgOV/+rS4BtRI7q8STeW
wGQLvAMrKv5RD0SzxCW8su/QVV/6oCqseYrSpb4VuSxgrOZnVZJV06VTZ0RaCISE
rgSrFdXUkTjBpT+/qeQRgGFBaMqfz/KeT5GekyUmtQUQwttW1zWaik6jwoRTxRPk
dKUBM71xcjgg1biRfeqYOsnNi9DCrp4+TNjk7X6Ap4QfYerBS+XRV+ChJCOaEQJC
nj7Q2E7szbs2doFH79iwtYrWSRu1SV+IBDCseJNLonAjTVR0X4Q1ZG7AYdaDCCse
1X5m7X9LfGTSjUn8FxHl2/bC3xCKHmhWx4ndWKz/GUOwz7cncO/pDMS6MRouRErk
6TbnE+MPWF3JyCysvtiycGjsPWoV4pliBgOnZP5DnZNN44MqOUxpiWTU6SRjkwGZ
zFPnlcEbCsffsHtXWfelP15AHY+qbkLeMJi5ggldH10DmgJRCQIOFvCAdcv7RPX3
PlkJk7wheB54cO8dvXMDHEbDz47FbO3dfxmrel+Ht7SvnUh+FklXZ5K9hU6u5/BD
E9hSvkTb6h6BGtvJ3Ju2A8DGTUmA0c7w11ksbagiZNivx0DBwWImwsB7tIbOTVB+
lRNeytYhV+FwSZBiTFZoxCiprkwLGZ7+BHZoG0WvcMCd6TqgP0/KfHS3gnj0Bl6B
VMcXUXQZJ1piZ9osgr8epyxjJpmUEuM+uhdCoMDUzhT5OHbpYWJ978n19VeVAOXV
sTel4wyC0tq4/NLfN099cbEoVAX78eNKWvQs+bIdDlwH5YTSqA/h9mvarzmCcxXH
6aKhy220RC34xyqLWxWncYiJegOmVFCvYAeJaxFZ88Ep2ya1tY5mhwQpXOq0OaAC
0cFhLrfxGH5wF4IH+V9EId8BRIKhLfLogB+RL/KY4nbnsuPfk3UTy5yzQZkcuXTw
q5igvB7lJRulKFAGhsy59Vs6gxl487P5BMLVzJFcSP7b8VhcgE0Rgfuyv4ViZI8b
jlPWPzVFVxykWjlV0m5sCzgPF5S50cwmoJIgtoT+PCGjLHba2WJsK9EnMQW7CEJs
rdlIqY5jwvUaqLVLHZ2FO5hhhz2Y6rNNypm8GB31tzEJBLQlrwBbg7KZDOT29PV5
HdcilaM4aqonu3+43PlAEaUziOBNRSZUC5SQEMt0qOnj+vsNUGTZIWhyHnRVQq87
mLoDkjyfWcgx9BWQxav9QEB1C8Wb/lX9lMBUX8sCUmyvPpJ/NYmEZleDObCtM3ts
0wLdj5mo45xx8s6W3gyV4pf5ReEWxdesrRSlPip/752/Z6w8ZSenc6scSwinZCCp
KelXoZ+OoW+Sm/2bFsCQ/GJVq0SRUYoxX+zxeEkxBxvleQFTWU9ZPN5dl4ysDR8K
ZlBxiNnbsCksHqrjksFoyANzaTsEzM4Gpd+RY432ssG42VUmERgVZTRFZ/nypsuu
EuCrt46szy45qVDFcLW7JjhtKmKJ1ZXo5tPK0FEUj66ZPEJ+aTvt5ZxMkZtz9oEK
udBf2J9VkpxEZyhZ7ErOtZw4ehjK+Y5c2bbYwo9QXaPodtt8oI+oGYubip4yFlpp
aizzFamkS78VDqvcC2W5fgZowYaAotYl7KR/jHccK3MwFNN5SdNtJTKUghr6TXRs
FEdUjDjm67yEgI7DV7pFvoa0enWwCoRa1pD4vXqPBQlw4Vo3MtSyaRhycaWsPCyK
rXAfZwhPi8JVDDTOy2DalTx/UDVgqvlaTz+loxHdmdzl53FnoAyYIuP5LXDTxt7M
HIttz91lh6OBfRo5XXCxnVDUsf3OPPwKgWzRJlpu+bB8JzAjbKVgeA8cf1/BYtQy
xdIrHPbfIJ+pfnjrq3mr8KXJP9ftYJ2YmFsb9UEc1FB43XxSBDwPD4CqfwFbH1E3
Kkwv5QDQe1ibanEuZdEC6Ug3Ddv+avgU7WhSbd71HPmahX4fFFjwt97DA+Qk1nSl
3E7qobfhlC/SsZzpuFSiVDnhWHyiQF0vpW1IEmBaS/bEbWUxGzDOpAoiAlKApx+J
YcLb9WC244Ag3DFALLWU5F/sjxljswqMh1dUoVX0Cs3CXsvY+G5FA2699qFtCe2g
tijbwbnIX04dGL7SOc80ckWbGeZXgGFyp2thNITcAxtzj8UBQkb/3duVtTuYPbWF
ACDS3nzqZDGdaMpryspKUQAeOKOCU97O050TQ78xV83yoT1KaQuKaIlQP0EeU9ua
U2vH6wHWH56NQKp2cb8i1VcIZDvsIGsOTMB8DkxFxOhJwRE4OLOgbfsxKMnxkP5V
BOlicP7BocgCgvMQXw7Hkt2AYvODUrcndOnmcy4fzdUoPMHGfCPJjMT36hVpFeDG
TVZn5MgfQGAvUaO+yw4OMRPW7Fl8vAFKcGyvJwCAJIYZIkNA6sHaVI10eM2byj2A
nWjg+WoU9J1R7bjwlHwA0ALErXiVea2GkBIBziofWY6MqUTsONRYKP+loJwh9lQq
bhbxz4ciPCXcYzy9oOgi80z1tYGVvIc/1ZwpCCLjJPDI8Jceinmt19XVtzS7Kwxj
HA7HFg2GBj6r+nBM9iVrUY00BjlUz5VOuNJ2VDwWet921A0x/JURM0tdUPS9ioAq
UbBzMgtIIcW7TNWU2uzdRVNxAS2AkbDagmxsdygTgSl4DaLZn1nNGAY5Jd6BY1O4
488ir/PiEprb+6BjYg6RTbPt2eopNhwDmIAKgsJ8PAlKKbZAYbN+G1jYJevVsDhQ
ReS95wPlYCBjnPV64+4hKZLZWuX4jth1msifvfdP0MKeh/36G962/ylMPi1grOog
GbdBwIEVAaI44+YEO4bcpgxGi28LPMTK1u9jl1Qtt932F92u3i1Q7zAQQ1pCjnoJ
GyVI+hH1vTzdOKQogvuK/WtEYHZ8oblTW6jb33WwXgx3+8HJu/KktInFq+7OdyoC
3LbWvh4ZmeIDetXWpeENKx+9rMjeORw8XHY3/RYmyv3EiQxSd1eJbbDIYfuVlzJL
yNxU4yoKOQe+870EiRlHt/L/qgReo71EUATH4ZUXy3teYxuvqTb8bcL5HYj2bhoQ
UpMuLnD4TtCpoe2rU8xPz87gdOXLBqO6aKVWDtoFr6Tl9Sr53FqgfUSbBtaunSMc
xi3ne6/qy5/+rPNuUan6p887KB4SRCp7vzN2roayMcNtOvl5Lus2yuqPn5F3gvTZ
0uxjuZpM39z363NumHFB91FgTGcJS44CZ6NdnC480bustqYD2r41Mb0w3+0zsMI0
aT80otkc6CdFPZQTfqmzdK779r4fCB7PS1DPPTofywMy9UtjDGG3LCS01COb4zvy
bCmO4eOa8NlFxvLI0nxZwlorigBF4soMfdwtWUlHndB3rpYEVsn8GPIHHGPWEIXO
yA66tX4TceVxsLw4otUkqJ86JLZMvgmcnJUhnxopb48CNVSVQlJ/2YYG/CY0v07s
7MPlZmPN2BH1ENHA9bdnVDjWmVaA5rQ3M2vEBIBnh3E5pdTMhRAflC4RYSpYpg2B
3j3nsnuJZ33twlUreK7/TSmVellw1tfMteGUti53py/LuQLtlySw6qK/k3lQMrPE
6ligG65mp7xR3QHdFVP7/e6+V1CcFhxQZqEZWh2ZvZ7NNJkY8jsuwsgHSmdo+cTv
i6E2akS1gv4uhQeEWXisqFr29B0mcmCAjmv1QzDQxk398qv/xDBD4PQv9Y5jZrp0
l5jYqGc9mOcEV5nSEMERLvpYV0U9jSFAFg92sDmHClfcei4X7XqYbXaqglM6QJms
K/3xoDbH0xjBLCRFrYJWrSwfO8mU/F8bDs/49b8nSWA4j61D91aTeFbYOZEZ7G6X
ZwSuy5wtvJFoNK+i02qXr8Ksa15+eSosHg937oaNHBw0wcNNrnncBbUVDehdxzgr
W7jBmG/7rHnTduuCxC9/DXKWvtkftYV7nJyXrYC7I8VpETR+cZTxDY4tXLaT+Kqr
MG5ijlgiOm+tqLnfaeg4ws06oI5Md656AL/f7sfxENjMdceT/BEfe62/F/jx+IQ7
+sUplVa9kHu+pDFBL8HfTHn12mxWad/aKDj+q8Pm1tO7+w7sVRHlSFGMLAKQCb6U
q4yz2BXt1OUWNYksLxdlEYWhqTk0kfCo06PDifDkqa9TRwRbo9wBtvrxf0DKu9+5
oobBkyn015A4kOC8zG110NEgjkjEy+0Smk0sGXISBySBoH/Tsqku72lAR4QSTP7R
KtlN7PqYKcnOlYLElEjTvM+yT3mNLvQ076sp3tpEjGDFfD/lCqeughg2vt572pKC
agDBRohA2YDpXX4hoyiuR9NS+gNTk5DFrU0S9BQEM+wBirgHNbxd/exm3UnEF3cd
a1+RAG7KbO/1Q9c+hhr1L8TX3IQT4qhto+lCPdVekqK39FcuaboFDf//cptfnT5H
opPAMokAwJkau8BEt0F5zUSykADcIECGrr0isO02328hHblcMOXkVaf0kww5lflr
SyszHI16bwaWjingAavjIoWuZogY/bFlT1pPe0iDwdV1izkypygUD8L8RttA89AU
AwcBqp5wvrV+hYDetJfBNgnN8dFD2Pv1QmR5PIFuCDlIe8dN7kJsayF0HfCAqM2H
STUhleLGMZjs6fVJzSS4dQdc0zeZqHAxJ1q0D1wAw+xNrF6/aX+hMhLacrABnLmf
W2Nc773VSGe7J1k1bXwGEuvHXpy/7linmd+uRWzqLrYIg1C0y2sw8Cq0ORFCUp6M
tyhKYkYOyom2dw2JpUmAIEWIB4X/PCzwCZn6vnfEYaBFonWCpkz6c6dbF1FbLx/Y
aY9HYuPX28x/vcduM32GOKgjWDViqQ5kT6z5mZJDeSiQDnSwj/NCzddFYZO+e3l/
AyIX4qUHM2ApzmQ73q9nUTef0eH7ptCAeBdn9d1VTJPURrNPDi4bdkHjNSadqBNn
wiqhgEH4w+E2Qfq6qhHjAdpVPP//3vU+HawQDbwcOExQ1W0e+qX5bYL5ZTdPZjRC
tNj4p8KX2xcsjzymBl8W0baZB7acuwBsmFZO6bMeF3L9MiB2A/9V6IBtpjgsk63r
9RHoMRKHT9yOOSEEZId9iDq5KkfhJw9rH9tEdnvMvt4LRdyQRhKivgWNfSSKsyCl
bZ+rZ2VfH7ZrEjYfKay+3iJ+khmcbdx1tpNi4etR1TW3RXZmCrVcJREryf7Sf4/o
GyTiOq5LQIXrAMogTYIY9M3KRlqPclSIsAuqGqmKIq1k4tOfmDybrNghnYqhHAeN
2HigSBjv09nCV0LvklcqsXi9/AuHKE3YPR2K/oSsah6gM+kvtWNbTI6E+DAcEn0/
r3IakVmSk2y+L2s96S74ZMoMQAMq049qOLcaVno+oqlovP3ae17RKEKjIuT+BcqV
qTA/5w/G3+/uz1Pies5Qa9AclehbWQtSqjayp5vP5Ccr6OsQPeY0OLkiih7jsF1j
+oGFSznnrnSypeSN/T3imfWHIKZAsVC6tAU1K5F++MlMIxe5Z65Zy3iIbsI12JWb
ar0RvxAsIpm4yVlZlhEOGJlOwXnJcr6iFSiJ6HcMq+kvLdUeymh3qZ0aYZGbO51Z
kPt/9rmNLmQhOmxXU2dl9weEFmPlg6PxiPk1DdWqA98jpbzXraIUTe0SZcRLEkIo
vKYvay4uWgWVt9+bJGEM6LL6SuqtKxGZY64w4mn0tgCIqaFUtTRgXhVCes0djZuQ
UUDj4PX3h7FCg5c9Q5AUFfIgYIoYY2cFZ+j7/tWefPSNfOsG+FIW+AeIjDc8/GoQ
I2R0QMIjimhEpUNqoNWAU3egc/biDYZNFfI06kc/0uBx4ReA5PzLOFYC4UXfsGmp
r7KoR73H+9d3tI0ebei9LZ+HbZcS+I7dLn+4CWOFsPdFtCr+XJJK4iYbD42KRFgP
zyOGW3dLbUazwLcntT8rH+4eWCEHWkIUgAvIdOUUrkQUDWaDe1tOL6MoaIa2TVya
SuEUjFetwA/EMd5oH6Oh+juIOhWcCRTCORstOmW54QkG0W52FxX+uOuXmD8ARwdW
LbaMVNPgFHrC/W2bVMJVZYghkEQFhT5zTRJuAj2SCEDSKUZCpk2Xa1PqhffJKC1u
CL5PjCrhQXpZp/eEiinlsgxIwwbck0elgD8y2HLpWkcaNgs4A+ipca3y4YvhrGF+
wmZDIpKNb7tgZ3R+Fm27pHPhfJQjyNYu6PFv6ZloccWbybIbOsUR/xVux8Vj/1Gs
KphCaLRxWfmJKgPxMxJttIxyj78E1P8xa0QYCpzqPq+h1NGHh5xONjDpWBCsedxv
NrgS8OauD/Ysi3BIie0fRXhcWydHjhoFDxJKRtqZIEf0/vlQL7mJyZc/x/2FZ+OC
rud2Lg6iCrreKBsU3SJZNiy+dlnSjjudycySROTRxnmfmro86U10VDRrQv4+KkKq
EGhtI2GmXPOUKCzfJnxnlaJNBPMq7kKJy61MbOmpSvhBUE+pkpCdZb8anp+EObk9
uVVxxlPOcnxM8wtG6InCgx08eX/mbrQkFOjgX0fAHpLEU8dp0LTTJ+fXmkDHXeeB
edy1rGJVejZj3d7UdUuor36HPt43F6pWr3ogtk1mi5Dwzi/6Euxdcb1UHgkGxBi/
Dj0mMFScta0Sgz4R+O0Gpt7eQInwKs6aQXwK9VnzV9M0+fI0nZqTOK62qiKCBO8u
t8KKoTn3M6nZgImjohqTQhEcZjejVkinY9m7kYJTj3SDD2f7AryaFUhnjKmQOlxK
SPMEy3Fxkoh5xpcaYzQ5y1Q2YcR02n/a0Fehie9VeUJy1dKatIbe/d1hX5XwmDfe
wJhunGIzBhLm4Dsq1pyx/G7RdtxszgpCNDJ652FCXPN4Xx4NHqlmjdicYP5WG7cr
ugW/yh/XRdayB/rsbGD5/DuuENkJWDJr2rrPh3Y6S57DrTkVtPmWXi8jchg9Mnz0
uUUZpAGIecq1ZVNy4Jb9I07LTgmISQUMFdYeiTTf/rvFnZC2BAgO3rQw/9XlIm7K
1p7819CTqllKOqvorn0B35yQxfBBy6plAxcNOy0IYBjKesZO2PRMLosvkFZy0GEj
xWH7rGJ6esYn+soJE4IT1ItnB+yHVBtzITUzoiyMN+QK5ZbRJjRTeYlrHV46H3xF
WJvSbsGMaqX4iWjwVqP6n+f2sJQ/hro0TWiEKL9gL3XXX7P4bSjr4f7pv3suc8VV
kCj02hXbeyPJf+VylsrkVjqwXgqNQJ1MdY5JfnK/WiWvlNOpn8sn2NcqUhTFymFj
5INAJ7SqZzr8YR+R7t4ywg/M/QzC0+0gtIg62iPq995WtQ8takS1/L/e0IKp7B50
Hh9a8AukSTOQmW30kfLMfQ6n8nsJrXRba//7dszL/o3joVvigozK39C1HJqy8ajj
KmIkI6CYgS0UPvsCgDY3o43EnC6pciJVboinDV9OcrxEdckmfZYjbRU9sd+5h5ml
qU82QD8jo7yZueEe1Ln3KyQx1XueC+5frdKUe7QMN3y6/sALA5mfsKS/T77esSF8
eNUVpH9otiEQWRTNPMkcHhW8LmwwPzkg5KuZpnmG8ng46EuDCuHrTrZRJRDXAVkB
94/jklPkqM3XkGEJL3lIK6SUQ43gDvlVkBj0Mhku8IoUEoHHb7VgDA/AUNL5ZwRF
b+Nuu7AhttHNtttXwLzodCQpy05XWu+5/Wwwqf6FIlV+/ymNERj9nGrPzVoo2Ku7
/XteDzCXpMRSw/pNqjz/07vrzxlCxnzNWrDr5leIk1pPFGRw7XDou63A7WV1bIOZ
iFZbd0nwLEiA3WijwYVrhcO/k35C6EAQFZOPn9dklZvZIpemAktdwIhZX7ycMbL4
29XY+PnEx/cWr4YlBYfTLTA/Ps/+7ARSHLGGQxixpilYkM7lqa38vImtHkU2bvq1
mmI41Lu/ZMD9jQkUP+AmB0ItdQVR5l1ufMq1PSU/2W1KXF2UX84IqlXMwHwvuajF
f6jTT1TouuC20OIpomz3b4FIsz9JqoVLhCc/s1tz2ylkWWTxySxuF/s0GbwG+84s
7/sDsmOF9juLg5oEvpLuGM8xBqIaDpGy6Me3ECYT7mRNVFwIH7tB/HSA+4hjFshh
y1teVani1CijO1z4RrMjNA+eFm1JD4fNrFBKKw06YejFK7iwmM7qKuQRm2j+Otzj
opmly0dgSUTEBBWkKuz5qQ2juhLtvjPSASvbmESS7zp6pPuhAgwoSv8H2tGduoxc
pj7Q1fZKgWfXhZM0ch8F0SWK5xZ1p5TDmgGOrgsPIw81AVMJJvJcddaHP+jtwVgo
wj0hlN1W7vlsc7Oa63qprjxyUGYycz6eqdrI49qpv+EQKPqJVES3hlojkfYu1MCE
xElzIQodX84ibqK+1QC8zykkTizsyj4pn0r4rdBDGtNSwQra9jUyxGxSVBW1SfbC
31npITEajVIQmD5UP5cm66EhqDzEThkceIglUShqophObMcBcUZZ9TeIuUoqEhNn
1FW+R0BN7/4l7/VQ1n9nFfnkVOlhDuTdVvqhk/SiPbcxTKR78BWvy+E8k/SuMWEp
Ti54rW6rePfEtGEpOdDXOddtyFCmaWL2KLNt5wobab3H+wHbjwZU5go1g5R8P5tq
9ci7ptrzeUCA2Hoj4BJRVnm6d1/ZSeXRsq3TRMFyBjnXF902U5WpRlovXGRYqKaS
PE7/NlsM0JVH8yrpVsxEfvnbzDVHYsPCDUNrau5Tgoqk11UEonzU1SXeXC9ESyIf
wtcjovLp3X8XY5nA3ba4BNvMSNQT2ERWk/LBSUZOdO4=
`protect END_PROTECTED
