`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9d9THY5PWeNFEQWBaPxPsFSZXW7cdUx0FMSXYow9A/UlDtf3Tc5PGjzM50wSxfll
5kqMjfXsyQf5aGpInE9T4jnkeQh9fJbJBRebsEh3cJZuKdrviXiqjvSuw2gkmFH1
WI3iawPtFhd29/P55xWZNorjUzPaWpfCHo/DYSarrDd8golVNOEf0Gj7bZaKJjAf
NyvM8ut3DXpqK6UnvEX+txEkgp1nrbyjchU5vWjiCJFGpuP3JrHqIH00d7z7TKqh
p+Omy/cTpgjgX/PE/6/ES8v0iyC3/DQ2lFg3KP/abnOk4P/xIDcUMrU2FMxIAT76
FqqO1oQeLSIDLH6cvtFkWGHrqmOSIR+dDo4xcj/8ol5nckfET6HONNgaLlxzpYRk
KsFAdJk3qbusQdx94Bb88B/Owk8zCnitn7Jy7b+3b+xNwZZf8uazX5RnpHYLfYD0
qVoYOlAf+8ARx51JCjzsV9vI3diQKOFbkIQt3CDIlaZO7adBGYfBLJ5ILOHK/yb2
A+pe6vTwkc9tYDMb/G6TDk7Mb6JebSHfmvcnYmPUnMdREvzxxXDU5drIeZnaV5Ht
ej1vUvmewKhzcAwj3W6lJgA74h419HSlukniBbg377750ttcX/s5n7XgnDSaIUpq
bE8tleKIJv78VRAV9P4hZpGSoFFxmDGSVZwT5Hhsf+kke8aUors9G2eRkOmG5cmj
tYCmH0KHEWQwERvvK/XR/90eey76H+8+OolK/qzCARX4x0Ew1IDURuOD3hAd0Ahm
KYSedm6XtzsS61yXqm9NQh250oyzeXuSOkMQ1kJG5gM+wL9dp9GjmrIk/WZbBrOL
CRjYrPqBeZq7TeT4JEsX0SV6mkp+XTQUw5rt+SQ8ZL8=
`protect END_PROTECTED
