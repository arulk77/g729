`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBujwH3cR5JskWn2T65wahO6jay0K6TLdpIehJSeZWuX
5lqidsm8Fzv3Rc8aulXfR34tyqSWwFojBWYVW7ypfsOx9JbgaokVCA/RE93+UcFr
eX7NyuQXSPdArHfqssv2ylxqXUKnM+Ddg+9UD32g0sILkPdAob5BhCNFh3gN6QUj
`protect END_PROTECTED
