`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42RUZs+vaasy4RpXPIfO4qrK1FmbQ3oe/vRAbWNzxDq7
BPRI7UIBsZZPWiu3HFdQCp1bLH8YODFv6sXYQ0UuyDBm3p43d3uYQlUlvbiUajWG
9LCkpwqHyDdZb7jjLy7Wop2bzEFp6MFZIQbB/pR5PPbE8sOmaOIeU09D8BWi4NVZ
rLqMrsp0VT0l4kfrMgS8cha69jqWwAPfADDXA/23505xsvjW53NZXnvwwsQvbl4x
40O4CGN4Q/88HVdxs5VN1ihnK6Nbv4AIhWO2GR/ifJT4lMj6zpq6lvt1r5ivrQk3
1AkICjKFKDIvqVJqYJBlRg==
`protect END_PROTECTED
