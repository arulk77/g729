`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu409DV3xjJXG6SAtprq2ZyDbrywUUHSC9N24Whgryeogd
abhngKYANM8csCT0Ytx9F1C6pNmkG931hgkXUw20GhNHodgH011BtYcYOM8qdpCd
ic7haGF1vq4d8zw/Gfh5A5spKPb0leOyMiamCY6uXdgQDB9ap7vkTatEfbHPI5Hz
Hrx9MzKqihl125ICLXOoEMMwlBgi8CAYhHWfVi9TWCr8LPfYXLH1uM6n/OlM8XP3
la56bTHj4aRYv27e+9zLIoUXlITi2En6ZLGkgWnYaIUsUkYKEFpStyHR3gSxk339
Kb9VXAYMUJllVFOoRfhz2Q==
`protect END_PROTECTED
