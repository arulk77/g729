`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
h9m3BkAcPsUutG4T7rvwvLdH0n9rcQrqR3ZUiBIw+wT4srrkQyxWEQNORSPq7VGY
gYM+jVG1MKXNZEiS/DeB8QiX2kJ9IruiflL/6OuuUn1171YhlU5lYxMEkFs+eNSx
JD+MreLgn9vr3RNZHuE3eb8kIZOLo2CC1zQSjCWKaWaxI188w7jOgsNK9i/9FiZD
jX87I4KU1vbs5KLPIcfci38NhNfPfXDCA7QTlUxhc5eELdGAmVwnQvVJQ9RN7BG5
/fDVCySSt0fCHaCcR+XW+8FRyGJ9PJEaMFPPFwdKZY5hhkIpl+JuGgwIZNK4J/5D
ojNHr1UDecxCvmqKOHuxtZn2E++5QlT4+DiGrxL7fNBdpOMXH0UgCYWgD91saaf9
FdhxG7IJvcmKa2JSjf7ZRvowFG1xL8DjpfrOLWQ5S4R7D/fliM6wtLichyu0Dc4g
mCrfcM8OS7KH0mBIN3GRB25bSX3PhARZLhwjvmUpzVAtkZ5WWzd2YZz0h5HRZ70o
soZ0Fmf0JZRqM5tWo7msIQ==
`protect END_PROTECTED
