`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLWRnGq9j4CTbFda1Wsd7J6EBU/fkB3k2DRQROhZCHlR
mdKEkIb1rgzJMrOfGBm2E4Gb6+1MZg7JdhQpQfgATLjleGMVFLMqKMDWwEGOn3QS
yqomi7fNDo4rGu0ZIIRVYWvtqNkMyndYR7t6PXRVP+xdkqM9JkQqaAes9Yow2QoG
XWdo5a8s6PqchMQcb3C9wvnYIsMgXdqlSfpG0bNsa42C2B+UbSD9HA+xivcedllK
ao13ECFThPsUvHoWiKZD+Esu19HBDHlh9fIN3Krda7tKRr7RSLE3/ZoGgOXGZcTN
ZrB0BOeO3ZLscNZR9kg3176e8MwvioTwVsYAadEFpPMxmAHFj7XnfA20ryd5iNog
a7b/xsHgZu2QwN0MfHFACLSZ/GvddKa5aWTDABAp/ih3FjmgxrHIw/fVu7qreN4L
23f9JmsHrQzdFGhYllkpCGxA9c+qbWJFdyeQGh1dvv8=
`protect END_PROTECTED
