`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAneeVwZ7QbvlEPJW9v43Ukw1c58GnCW53XHTOPtvqZH
kqcAxgt1+KQlpwKYkr7MZP4zufJEIIOpDXNPksiVjdcTM9Y1XXyKfPQIKhcO1/Ft
TAtBVqG8OAcUyKj4iddxtxpJfk/keYJuB8f13i8qNjZAq7VB+vNZGGM8SrW1pTXr
PYO75KCBHSXEw1fvaDg7TXPw2rYYfaj4CZHtGHyjeK1Fq4Su2zKg8Q3uoJNFUX1e
fhs8L0incH8C42OKDqZnYEeSYTUikw5ZNreyybeNy9FkHCUp52g/dC8wQkISAet8
fgBtoxnT10rRQwH/gnmKLXBCOi1OrCreGJD7yy7VtuBtfsnrkT6bgYt6GRsLKaMC
wm4Z4MU8Zn74jLPMU2fOrE9MlNrTjNih2hXMt0WYv091WIlXL063WcxR2GNRDMwx
Rdabu7oG65gTDdRi0vhrfySnG0W6goix8Lgz7PRsA82eNXxc207PNAJO6xDLZhvg
`protect END_PROTECTED
