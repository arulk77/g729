`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIi+XgmC/FgckM79ZZqSBGKHKGLFGWPplH0YBW5pLN/R
q05RTQvPiSc3ksbEnOgWU3bKF7U40hf+gsNWdJPtYrVCSZtmZKKBkalMs7YUSJtb
vsUs0ZY4/4pbaE4h7odffYrF3iALUwlh4ePQCxqsMU4B/LNjEOZ9OPRXTGgN+dV3
7fVQZI/mezjPXbnkTUaMZ3QqRIzLZTOEln1vJGd5AedtfCNsdr58yTeBENeHpd+l
RFQGy/dZirXv59lLN7st8SVWR/WFFwTrpgo3DUGbiYoxt3KaM2XZldmR4CyKE5j8
+68Vm3qMZqCTETeZUpkMHEY1VQ/e3ZEEBMjmNaG7RLZBCsozTjfq+IV3taSNdnkM
25PqZr0CFD8cnfxh4dIlU0PjjCCyM/dxd/qw7OwICDsNckWxV9Y2JB85c7KYvtRc
RMjp6Ogg2u4w84z2F8LGwxtcchu98af8gQeik7FNh2bVvMdk0X1JagTUmWQ+VDOP
`protect END_PROTECTED
