`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOrV6LVGLqq94yc64XUB2Sz8bxJaNlaNMjHWJYOmjU1V
t4yoPcb47/4WW/9jVaod2a8LFTwjcaScMe+6BdTf6JN03z4XaGj9KFmbmBMNk0ro
MLvz/AENJecMRUNtC1zk+m62Ox+4TlWxadxSQ6uGj340XN6+INIJhUzQkDiyigu1
68gEURMCc288OzNgatlbFs8jEUrPEEUqZqBYXtIit9VgFiavJ0YDNffO3cLEVF0Q
+Eb6/SCOretfZIYQ6A3ApUzk7+/8SCAuQLlSK6prSyBVeI6tFfjMdkgPChttjix2
UIt2DHmAkT62b45fKTQaMljccwfzGNxrkVsFGuutZOBn13ILUY+ZckMk8Xka9y5a
7yuGo0FCsXB+gizCTD3ekHMGmjD2XTXs1giurqIA9F1cVMXHxrUFktlqEHmDdlZV
mT2Wj+Ej3v5hxW4sd4TTnZmGWyBtOPicFSUx8eiuRuh1qxlqB/ItpzFbK0eucg+9
DLYjk+oY3v09rZ0hLa1b/St1Tm8Ab6O2y/S32YmuMQYheeKewSUWYpEddoFV0Y/I
XGHIG8XAPSAhBKUM1ONZ3wq7JmG4GvSAjrEzKjkVs84DXS/0alVWeX628iYlXhy9
wDlOSVY1zNebB+aleM7Vllpk6fJaCpC7Ptb7lFrtI/FdOM4FRX/meKACTi2rveCX
etESDbOj3ZOojsekm8sbnbANHuckBal+vE4Qi7Q+6gbtd0vmsm4O2ShJzB1MqhIO
BRYno1ImHDcx0h7EcOzU1t63MepIz4WnAUpOTtmzVFx2nC/JpJ4JpeEPtySK9++I
WTUKXtKjnYF113mrBzC1H4mBxnLUWVcc6stUKrIG7/E=
`protect END_PROTECTED
