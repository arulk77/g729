`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/+JhDQSGZgvcBXGxjkjB/3v/oZZ9uJCVEzkPq5t/ALg
2BpmSIQIvv2VGeWkLcxfYygbaAGkkIrVjDaA7xIyef4GQlw8qtP/BaKIOvwrf0WK
mId1VAJjTdUKO2eDlAA8dZql/U0Mvvn+19uSovY3Qd+yl8ws7uvRuP/mSrGFfiI3
WiYdwO5LZSMDdZlLS2JSMNrmIfs2d/zs4ndZhfDb1Oo9pvK+mqDoBR9cEX8nRjTO
P3LwvxkSACHbAGdcGa/YVYOP+Myk8AJw3ijYYYBBiv5LsUDl0xqRYSxUsuMoKXIt
PTilVLpS+4F7hIbVnzElHw==
`protect END_PROTECTED
