`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNZw+TPgeLxkH9imxmuYu7SFMrrnkaTIxqdnT/v5JcJN
V7vLUaB69NLCV+gy/g+fRMqPx1kH2R7W7mKUwWQmatjBOWZAelH54UimqwGkAU1s
wXlG72aqR30adZlpRU1FUIdxxXuqD+HHeI+5+4t4ETo296RJFQUe5VV5Slho5557
APvzogEDY+qT8VCk6ghe9lVCRCtFNnBCqXPLyxqJdCqYwF6S5pU+sM0P9HoOp9Ay
LKN2DcxQwSVxOwOMKfIjQp/TOYoyRtfHdoymR/x7jPbtmxzXV4me6VKNgiCJ2Cze
TI16DQEUWfJ15pw763+dQ9DwOA75UHvJASAFRc8AoPGubXpIX9r8C/8p59oMEruE
vCeb1vRApyfWCQ4Eqaz0hLI8XDvDcewsnCIQNo0J4CSrcpeatoRuoUAk+vq9aOdh
WqXn1JRpauFWf/PNPVYb4nO9+vZCywsu5u3FkG1Bxq2H1Z/Lh+YrKvOc8k6AiM8b
OCCiXqGq0njixEpB1b67YpexBmGP98p0a/Iror28NFKIkH2nWGUfpEoBAq+1/2LS
ZvfdjEn4zmMl+LGSQcVo/6MZib/3R+M9Li76nKG1WxOyWQOCajVQf98ro4ERxy66
+rBZErseJi1Fz6nZOjLF/ctEnknV5Prp0qsaddv0Mjpu/hEWyMvBHiKdTi9ED1DC
hUNZRzQAFlx3XMrgFNZCy5sXLfYA5r+AmghuFdY3NY0BA+frWOuxtfS5ONhZcmhp
lWFuq1Gplg0MkwnhiZ4SEhsZA4Q/eoDjwRLHoCQLGkKvVwWt+idexfMBg7yHjeqM
Ik8lpurjiyAOw744D/OMptgIJf1n5BPhfx1PQFuv3tk=
`protect END_PROTECTED
