`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
I8crr5hz+cmuvBqSF1J/d2WcBMy27g4nrhRlhqCmvIE7eh8GJe322qHUePWz0mq0
huwePy0pJa/KEnp/wIoN6ad7cKFN32lYECdGbqk7fZn0ipkdECXvHEm0Xcd48Jls
fU86TizN4j8OiZWNdVkBBQIG3jw3N7Di6b34YTEzvYi5FzRXrxy8HlHzsk94ztf8
bHQMNLI7IPxeXoFLKqbHdQs7c7UmILC3JVTmNtQR0rWkyZLig1WDOww3GeXNyJAD
fLK+SZIpZwu1h8nTBE1qc03M08GdY/nFXr4wIFnqYZeDTyf0RGpoYm/0clfiOTWn
j/yMcHMECJG74GR9fVkZ+3Ubp48ro+czANBeBmxZU/0=
`protect END_PROTECTED
