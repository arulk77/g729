`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGFexcibhT76gaH4ge2C5UzwkGLWTirrtRvay7jGbG71
XYeIDOCDTq0OtaGSoNOWz9EoB+eCrwgMTxLe/F0U6YeFHnaZWVg1WO9eiRYXtA1b
37kwSNdgJKvv+MesFRmaaNn4IHxo1x4xz9MHPSOpj6Za7BR/M0tR+UM6atWbKnei
14+Qw49awUyMQy2hXKg53rjfR3b2fT/fi+LP+8DMTcKrDCy1c6/r1znzNRgdYQcC
nf8zDL3fs7HxweHt92NtbOxJgwhNA4H4V7SI63amsETVVyChHqESJuKJkUaEwCvY
UA3KJKF3buDi0zdNFuGuAXoXGKDg/GKwrFXCs9J66TTMDSe/mprr1OwsuYiabBuS
WxIL5ic+OPMGjUlnZ8vGXmB2obTcYxrl5am9wMKkthWPqfWNi5t0Wz8l/BgQtPl1
+9Vy2ZKqKHBc4rNjKm9L0Gn3a4n5BasqgE3OZEG01q1S3zpfOPQBY+aAbOOTAL4e
B3NvHm+s+pagQ8JBZJTjrPzUfPv9ti9BtmtcGxmNHxorOt6SlFncmsPaMoKCLe9A
r4m6UTMNsMpXuUbugpqYjg==
`protect END_PROTECTED
