`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePbAlwJ1pGJsx2rNkV9LxVVyQ0G6WRIJEqtCMJMQBRrp
01s1IAZI7/xqOp3JVeuW2EuaLntmgQNwX1FEI/1CM80h3gSySs5i/SM/XBKD/jDA
EdCknH/rHAXzxKbz4BkcOOsKMo+8xrinYy2CM/ic+4GSRfaAQj3YqP396to4Ruvm
PSEHkiDdpQGRO9TN8p7IPnkeR/y276scotRNI0AIlgxDDsYRrF0a2fvTRIJzotgv
`protect END_PROTECTED
