`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL80Q4wWgx7IcUyuJ5gKhTsfaON71zG+pTq4vtheTzbco1
eo1CJBXrHQQ684MO8lJlPDt6pBzFG++XW0ay8RfM2Ty/NB1ajCeWophxZCQQq9v+
1vB1JGjxGrjXJQxapgLovz9c0HTHw1/8l6poHBC4qvEnEoKZR00SXqyGFTsmhp7X
x2umx5jinuFi/R9cjjLFuwB6RQhQfksuyEkIypHCK1LOtIvsgNvEx6Rc3DAi3EZE
Jij5Qlg4a1vrvquLGjX3aj19pdszC1jLdxdC1Sw9S7Lg6/Iqqa5Bx9BLMj9QDLlM
yvzf8DmDOQDluIZiwESKIS/d9dcesl6KyoOuCGpcDh+8tlUCA+Ys379o1vt1ywEs
lRhEtO6Fh98d0Yzl7+lQiQ==
`protect END_PROTECTED
