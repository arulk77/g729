`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Rdf6imuG5v1SQCgunE28r12p1pisiY3LXsY02/l0yJAMJ1CXCu3rJNg3lcvDwjN/
8t73fosn5iNTQJtEYRVWiw5xz6d2XovgciyrlotDfNZ4ieXSkwO3V83eAaQsywLH
zR+r8kxDfiDZU89o+riHP243RasoZX9lZ6y/9vfxdErhk2PJlGDxU0+OF4MpUeq8
YPGpDMLKa9aKdJtERvu+FjYNGyytLDHDvZcZIElIaZgVEcAmSUoNX6G0JwrY9WFp
EvmU1XY4Txnu1wH/m5LvgbwFY0h/UuuaXcqlcGMHWGPRIwyCH5TxYtjAtcm4g37p
`protect END_PROTECTED
