`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
l8VZkFYXujvziiOg9ll94py+ehq30aegARgdEQpX9xVqZLOws9Fq7kEsRHnQDS2b
lOEqvztEOAFcMzR1Ju2BllCB0zeODLo+UFAi9N1GwpyM4/k1Ifc1deBOkLSCuo5E
JH+lZJjJo8r7X1ZXgDw/WXlB70AIiF8t/ftE3RBE4RTtM5+HTWdmD2AkK+7AHDeN
oPDEde9llctoSn+JLYn8NIbziD0wk7puOCbzC5JfuKhaNJPeYVtvMo8bSRgh0fpH
WBmlkYLmWuWb12iKGc8J57KdGBYYfw7RdQWlicy7B4d+jBTP1GFm1/IPdiJgJYN/
xXH/0Nijk4zB/edgSPTCkBKmqE5nBvogLQxx0u2KlzU=
`protect END_PROTECTED
