`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/HkL6yazHelBJmv6AmRMQkz11vfhj9Mp/4pPZV5b7ks
HPc+G5OXDLMVWM/lP9JN0AG1W1ypIzwXQWhV81ACcWMNWXFk8QIW2tnQt9Dzp6Eb
KGxrNNf+TfxhQgNUze9U0g+Dyh8blBXpRd3OG3u3hBvV0M06lKKGA6oadL/DNMjB
EF3/3XGjmWT/ejxpesr8I+3WkYzYtLplAUXZ5tJyiAEddHJI4yJW5y5qDD41QsNd
xvZjt+U1JvKMhlEH6DPjSC6o1UCw0FGsngj+V1GxrnHOqKjx1qPsrqSqwxQnQL9b
flK69NjlvhNBuRY4MSD7Jr6/dESQOpDUXCzIUzVspXHbojUawNgClDthGthXKSqv
Ga1VC3Tml+8/AHheinLBNA==
`protect END_PROTECTED
