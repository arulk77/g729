`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIg3sHOrZqQWZJjw6lR4XBNeNos6rV3eGof3g4ZdC9Pi
JQrd3LrB5WdP1lRlarp1lLCnX9t/Ea0mFhJdVr28QIMzqi7mRgVWCCB1at19OABP
B3QBjby/agx0zmNmvVG7L18Z/tSR9NwRfHelQz76JBba9P2AC2erfjLD7dPT1qyY
KyI/suDWHrNFoJfZCuTi8sajpWikXcalSz8FaDHMOSAi8MWLDnI69+ro4VkhZDjf
RmEFr0tINunrM4Ns8yJglivxW8mCFc/Jhu1S+PpTLzzBQCgskKsY41azSVCCviTS
Of3p5v9qhpblCJicenQDmO6pI+vp/kduKFVp4Q50b7ZKc7xMf4B6RwGDqApXaLxT
wcOh93qCRTH4FriAnBkDICh7/bDpEUGuru4lsH1+HtiNzQ0NFT9D0M84Q0CgXsis
`protect END_PROTECTED
