`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGzM/lR/eVCEhEwFNTxeBF1pw9glYN5QS8JkKLzBrvoT
j1Qetudnu5BXD1RXNHW5XCDRlgqRPi9O0PXU0r//VO3j4qN8VHFnbSgYXflaACw0
LduZ7kovsOxFTRJj6PAHLhMCqWFLgADWgB+C3rlfgqMn30q4QFFUyjox05pmoKh3
51W4KOkLioHWdgmYqE6dsFyCwFMjtn55B5pgbn4qf9AzR4JMXU44y2DzU2dPrDmv
9+gvNx9dcQjzIL5Qo5ePj72+aqcZYV1R3rEBHLzD5kgfLGXu9kxDDQ9cNfr+stOh
z4VblMNZT3IbX+LA6GPVCwscJyiLMA5NMvQVeTYrim2WpePE+ichfPP4tYvX9GLL
QCVwsMgPs6v4AA11Q5b/mQ==
`protect END_PROTECTED
