`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yb8+0WfvupuGsZ2vIOkvu2j13IT3Yj2YDBbf/guZ+T2
J3QfebFp4wYHPRADrJR1yH+b4cVqm4XifwC8iw+iogikAyhd7nkwnqJaX0oOU6EF
sGvq/fi0XOTPM7AXIxy9BxKgp/H4Y+ZS9gZghCbmtG09uAPGgWVQwiHTSQ7CuRHA
rPl2vv7ndbid+ieETe8fuDNV0Atwb/y5vCTQbv5V21GWsPCxXEDdS9I5w7gyD+n3
XrMVSvuezGE4QSgibUf9A+KNuiP0FxZomUZgYydZplE=
`protect END_PROTECTED
