`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3ON6twM0bRyFDJLDX3TyeoEIkFO7pm53qtdW2vMVc45ZFT6QGZDZTnmyCt6YDsBW
3ZWdnoNV33m+EQcEqqqfBKAzrczqZtmII6m0C2U4fd8zaHSaVKpaodWfQ4EREMcF
j6LuR8PFaAi9TsaZQCBTXcqtnS5DYzLhRFhG64vKc8BpjxDEgpj4CdZ8A7UEpPVq
X21GXws4zMITskURwmcAGA==
`protect END_PROTECTED
