`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBCB/CxDdxyUdvVzoGu1cJN9xM8WXw9bSeWCXbN7i3+E
F0HDZ3aZVRbAUl450VV2trXsnHfDgPvDSp9IwWjUOKZL1noGdN1yIF8DjkcMfTYY
/UnwSHXHw/plbNbyUguY5ePLvQQU3VnPo/nGOkV4jeregwHt3DnjviR3cE1EUEYD
7YMpYniu+/riY+BOCqN5w912iCWEcYyi1E1+QkafGGWzRB3ztIXuiwCYtR9x3PVb
H1oMZdhlF41LuP2TP1Y8BgmuSfEbeZr6lCKmrn9A22PWTJDSyLFSrRfTL6CeFZR5
`protect END_PROTECTED
