`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSG2SoKNUNxS5BgCicjkuQWG+dc/MjquLwNd70h8EZD/N
UUgdlAKyqcDbPs5Ff5RcjepXAvCAKkI3EejiGYHSBoQ7+NJEsc5BU0NmTJDYRgqi
uwDqSmxagfV+XyPYGj9+ifOKrMsR9uRvWas+MVC9n3p/mpbt/Lh8h77VEXW+xdXi
YJAVNKplRgyiBUxkf9xbUsqWT1rk2J/CrSI0VKA3kURihuwTr41ukBiLxCkGtr3m
lT1x0YCNQklRjcyWQYBu/HVhD86qDXbYC6pwqxKVajpoyJcuv1MnM7fZrgrkp9Qb
tdhlNYbC/5wvuHsgWHwYJYUK86HlJxCev/eBZfE8zJ/y2vncBNbNC6gyVin8ZdhB
WnrB2CSCmAnktClKVgG/nX21Xfc/lEnDIz6l/FIc1fKO4kpETINLTJE0A5jOC0ts
oalh3fESmg4pMTwdrjDaJJsJJ/w5spidj86TV+6d1uk=
`protect END_PROTECTED
