`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDCdN72pRsuHgoAlVbFalktrU2tuZSH2nVBH4tNfl0WR
cv5pM68nJ6ZaVb39qlAAxoiiB1CvfsVh1k98PZnr+baL4ZzzkuDdXahZjbdbZ/+J
mn8UE5FRUKJJTbPs8128aXj2RtoubmOUtORSCZ1eejgHO4M8s4llHtSJxcVl5i54
JRwcHomvevqfMZ1+cNVb1tB3JmxSR/W43UptvFeI48FwegHMV01slMtCxDHK2cdk
3PLLPkZJl5X0+Uo0/gg8JwJ8Kh6d1mF1mZumGhIIhWtg9IEyj4PtFbG2yncfy1By
yefuzDL7+hYCNjR3Usp6N0NsklofKpsf6A1UteyZuyc0WplHRYl72o8TwrKvvzGG
0MWEjUMUj1NWK61SH69Te5j/gAm7zpmIUmAWsDgJGUSaETrLxi7tFBSUPjD8cyb8
CSLpH4SfqZRkHvVbCu1hHkzAhikdUVnz5C5lJmVEe30wQjbYWrERuazGsHfcGU+s
tJThdBo1pKzJMaJ3lVbQesrp7T8BOf3ZG++jRhvrNkpmY7odS+VesIlKL/TTK/5T
`protect END_PROTECTED
