`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJcXXt5NkRTXkePiwOw1WC9eCJhaG9/82cRkxCTMI2yJ
BmFjCoi7aVM6NB8TTwM1Fywx7/zBj4rbYj84BdeVFS8qhROFzVig3j6ucTjj92Bl
BxiMAWh9dnspi5vgKemTPaQWPCtlAHzpfWyRwoDStO18TxT6M5a4nOsWDnfdsRlM
kb5qExF/X7LiArRfXODEex3eCnDLWLYuJ7RRmKMKZR5qEgHvLABlQBbId7ls/HIf
`protect END_PROTECTED
