`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIKqS9lFtf2wHzUv2dMmjEtx2fejHQj+pkBpwB8+TbLk
4lbNSivfxz3LDHmA3h7cHf8kIjzkpP3i7ODd18KhNx0ji2VAwcuFh4cjZgTKsiEa
ELs8dBGXcCeBjnxvXxUf1avTmvbJAjRDAE6J2LKXyAMH3qCGJHXPmAxTbEPdoXmQ
8hZkrbMDfWW9Xu5DDWB/OQPmkqS4QYAjMByjdxSO2o9crgymNVd6/z/Xo5gWTzXb
r8oevKh5b0UIEJ627bgKCVWC1WlCIxVf98Xp2sVmZ+taFomR07BIwptgEs0qs/zg
Cm+BFLGC5CeTDETFrRDeXlPaTnggAOnkupYMH1sVQ+0vt7Jb8MvRreWbcqwSSH6L
F+eTzAbFU544q43P8b0GJK6bsYnrijOpUQZecd4wxwCCEizg8lV9TfSS/dPh3hE2
shhlMdyKy11Qg4Yalubqpe2uC3DFKLf6aJRRwclpWQysoJ45HDJ7QBJZvg01GzoX
gKjUiTUCnR4NuJfmbpCPDD3WRKlYKWSZhT1ZA1C9WLW0j3Pg21V2PRWUTX+ItR8c
dGKm1ck7XRBpwmFNlAM5HdSegqBF7/a6PU1QGcnVSaJnseIMOd+y3Wm5AiZkGqup
fsXDd3kGydcsJvoJW79bbBHHpbl26T0MoYsuF2ts5+kgxpmzlsXHBB2UrjsPPlZl
tYgbIje4EE82Ou0SrTy00G6AAJUaUKCAsphTXMTnR1Zd4ML5w9g5pbKGWxi5ZdfL
HeFKhzdYNMYXptLiUMIrJJ4Oz5drsq5GyI4YHkwz5RMcSMutZs3QpVzIRS/t4TTh
6uc18tiSxkB35Q6JrV64+Il5+Gq9Vlizj6eQsdXyLrI=
`protect END_PROTECTED
