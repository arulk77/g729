`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48gsC5B5NIofZ4JDtogfoWa5hik7wbOQplMZ7kZuw2pq
MOo7daWj3xjtMQkiytG5RAcO++VeLqItjoTniXcvbixpSfk9MySzC/xpyO51bwg0
4YjHc6AtgjI+LPoIfk1mUAFWVCOcQPUeC7z6BJdnY5sAwu6vbSk9Abn1e3zwr693
q6qXLmJHlDZvwYzg0r1hve+ZAzFHX+3RTEzCl9BmYtKgurSGGYqpXDbkkECaZ7Za
dsxm9rCStpXEJeI/5vDsnq+Hb64L/rlNKIZXmpzUquIw1OfAulcIwQN4Jlpgjuip
jdxx8DVSpDKZzPsk2vcFfQ==
`protect END_PROTECTED
