`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePAP0F35ikE5YIV41hpa5Ms5FnhO34/6GOXjOzgzUP7A
G5IxnFECc6ROu4vbYtggmG2dWmKTRXlXmzc+bJDkdd6oA/Yj7/MbijnwF3UwtOrW
+vfbyPFrh2uJPDxLcmazc7jdVyI/VhE6HhHkxeRfnad58Eca8LWn7jdbrB2o6Jk1
8Amys7JpMLvTdc1aYON+Ezhcy1bLv5PO1H8woNlawr/YHMy+NsMTmcm0u58xC5m4
`protect END_PROTECTED
