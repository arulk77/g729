`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOklgupy4oUna4gfaccebQ2Lq7nmez+zD3BRI3H3PrbW
tXOgc8VMNII4oIWAV8nuQShaRIRdpAcPALXgI5AxEU93FKyLEeyZok4sjaIx7inO
h9UPgaR7w3PBfeTtPtwumIPk9IKMO56If0Evx1LUl5xyJQtXuNbV1zogrcQRqEpF
2pduFkTZuy78VjDOkpIik3EPeU10W4yA1X3MsFc4XYdegCEUWbIps9uI8ySe4LcZ
`protect END_PROTECTED
