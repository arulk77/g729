`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Fic3ua99JSXQEWrTTLOI8TIPQxyOEYUmrhka6kn79YvOD2jUxjHR1TT2mbnxW4Ch
7I7OHbsilwGAkoFUdNag4rrYJRFJzvcPC67lTM9/UWXZOUYBF/qm7AdAOpBvqWH4
eVf0j9l5ly1FyLtqWHnAA2LpnEFHq7duf7DyywyODQmU0XXgHWYDtPJEt8+FRlht
BVcT5H6nzYJWrF+0s+jaYFV5uHdX/VkLJiOG6vzKR7wGAyfT+J0Fv+oElfVhLam9
juE4wp8MUBtJcsbI+hx/CopjwLGDUFXWIbJ8djM5e5vhWi1UMOTvSWBvyG94TpB6
FOnWXpw0mR2NhlfAqK7Y/T54+klBcbtK6HOCbUTxaxeN861v/iMV0qFPFp8KJJrg
5HLcAO7/5a6voWv+mz9rUYCjuS1ruJORXhbIGvQHcSZ9UXXyvX71ov5u4Rk4kZXp
3EodMDzWu+l5mLBpjj0t5VgpK4J4zXzunPo3ihU2GZ2JAsxql6bZcVrlgxjnNSyM
bx7YzutXEaBuR73u3uguu1PnXcldzgOlYEIIPa1aeqEaF4pvcQ5he7lr0KJ9fLFN
98uJPehSrim15Z0xYRm6Sg==
`protect END_PROTECTED
