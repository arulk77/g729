`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1K3ew0Og95u4L+4aac8p8ixVgOQHyPzJsaiX0IcRGdDSAQU5IxAQmEZ1LnyVSm9z
I8V4Rl6ZmanzV8u5LEQjLlttfUqvYce41eS84MuCdn+Kq4oRELkClPjDyB2x8Kqx
U1th2puaVpMi9F1z3R2aT6mVdIDu1LtQoJV5GQh8U8ka4ivcS5vNVEDEUa7BIDlu
qepRNbp//9kO7N57B6EhiZZKYtnqgGE7R1sQCnAWPjbrMH80E47mDSzeR2ilib+C
U+MpONPD0xQNg7cUaAjM9EGoBa2C2QfvlmDXVaRrfms+tx17YlMAEXT7VAgtE5Fs
S6FX18RNvS5+O5pcXzimJiaZddmKczuUxFgDM4SChasrSlgJMGMpIzBR+Puc+tpH
YjeY1760UVKyye7+ItEXlQ==
`protect END_PROTECTED
