`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43I57zj52sotaQyOsFqcgr2OfUH6LSwGRqvq2Jr73VUq
L2zVpPG7cz0Z3AfIuPvPNtXEPXsXhYeDXmpX2wB2FMb9rjkf+VKeOKYzadbcRIL3
E1KbUzFm6kz8QpNEGVxHKKPovWDpzk3kM9gM+7o3bt1hPGCy6EKcO6QOfmoeEH3g
bMzEUhimYMFvFSPxKYKlxz7V70fH4W2UwSVaE/N6ofE=
`protect END_PROTECTED
