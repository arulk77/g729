`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL6KvNlAgrVyOaHvu0d+xkRPM5UStmbe4gKcXaPwfiR7
+6DAbP+d9+/QQVkzoCgoDERrXEKsjUCiXIBQjmOiumTB3L8IJROTg1wtKbsd/R1s
2FrDaiklC2frwNEyqMKFSdV6gHeA4qBrYZAzw4p5e8xQPINlplGC1BVYopt7FL3Z
O16P5XryKrD7MbM4lbyt02yEurNFpCoQaYPptOKkPuuNEieTvd/SMb5AZtNHjc3/
S44LJfwslVH0+zJLMx1JDh34OFvo/oznBtroyepclmiOKZAB4KEIf+6i21Z0z4GX
Z6pb2jz+2cdE6bX5kZd0v178UXOG8qqBX0WKxkzrVMgWo4hKDE/vaNUyOGF2B2tc
zjPeUeC0i63FNqt251d/H5KrQtJQCso81zOfUCARTihdKGOdHGrpWgqowFF6cD5t
rhiBJo1GBOt/Doegxpe57a/EsFyHdKYwef+q0WqusUFDHj50PRsEa9S/j9qTn1Bq
+pZUtNh5Hl2O27zWI4qN+m35kYbwUQm58UOa636vpR+MbAjF/OyudfS4IQ2blPfJ
`protect END_PROTECTED
