`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGHp/veHeGCUGsOHgoej6nAE6VpkAZMjsGTFDg060vvY
m0u1PsM153qwXFPzTRIpyYx4LSX5SYHUnGU4/gd1/0Ny/CVWO6rUhgupl+cC5p5h
2ZsbC2EsHcy37wrV1m9JjkIIDEk0Ub8OTg8PmdPDWlVlHcZWY6yyCIvu2zQm2/Di
2nvu7nAakkWQq2P1Zsog8F850iqGvmCGBCqbJaYiIq833KfDn1LzFgo3R6f78lnY
hagmJ70Z01myTccQKNBqWgsqR+cuvio7rf8VvbnpdvadBpEFgiE0o96IGVtoUIdq
iZtC023oZdC7G65cW9FUbVNQnb6vUmTrbQ+qbBpQslVc6RB9RiDxF399E1wePLvx
DmtW6md+l93EUuvYRB6V+N1RzG2mmg0/wlJecm8Jb+O9HfF3TNDFY3reGGuqxpGs
L7z67R+lryVJOxSHTGbkJRh/baFArTXffthRg9tXZQTXisVyWYvibeHCrqRmwCj9
3PeEqhxCgReGmyVO4+u0Oz6ozDJOb4rLFRHPPwf+tc9rsJn/a+ikFUxIaQTQQ4eK
Oe4AON4sIkObJsMiZfejBRLB1affq9as/cg8jjqvyaY=
`protect END_PROTECTED
