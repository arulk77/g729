`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3FVIluJlf9kYhIRAvK6asClcCexcxMiqeC7RTpqrT7U
0Spymq+biciw6uWAvYiTEwHaO0I3Ep1DRVHN0NFH2+dlhNrndtlCY/A99yPVTA/X
nw18dV0AcNEBIyrF9q5YRyRM1dkm22m+Ki67lkfNeDPXCvje6xqfDgkp4BG4ClO9
aTTMpD74R+2bokkOF0m7zPga5Bt2vxiJGB4KWnFvGVKQ+yCCwB9Yh1uB6Mtt1yEI
H6b6buB+SSmCkG6TXSexnMcpSnkquO9AQ+BMtqZVfYMkKVb8fREo/nCZY5I/bhBY
ydeqSrSOQ0qfBLRBK6nHrAvyVBNNaTyoLXzRBsRA8Gy+tu05A8jpTYlTWA5bwcwo
efa4e8xZ5PBRTaydVOA/LBl9hwHIsmTZUV5Ktw/WhcxxW0ng5PrQGWvsiQgvKH23
VJuQ8tUjUWRaXtBxPjBzxV4J0BNOnj/UUS5YnJoNwY41/hqSZROIV3r8dRfLuaXi
0gvUFnD9P7LInn/fgwfVHRshu+y0BGm4K6r9biTXbrajWWMo2HqogpQY+VTCOjuV
T7QeZh243Ius+7qgFgIMJ10KbBLSTsBvH6kei7wvugxTIpiWa1WuBQ9LF6vnyXNG
KqYzWmtbBD/S9h0qCcgV6zgaBO/X22PCHPtvMqBgt9i6CJ3hoKgPWJKAAioh2YEA
M24S8djzNy8/uqPc9s9zbbvbi2x2nSxvgnPWHWfEXSjf1s2ZBOB1GwM0+zjJHTBj
QTjY/5lNbxCXH0u9e5NRLmf/LHG6eeW0iCAft6K+KbqkmPdyfyBKod2bBoBEEDH/
n4a0mKCPeTxm5IO1K33W0Pnzs31k6wEy+WZdHt0zuc8TfpIovMG/jHp/kb+UBoEb
kNLjG30zTUk81zxh+ZgVlDq/IrTmCRtet+LdFKUsVydNTilhDPGEoLtSdnMaIiw8
eF6/FSx+D95Sosc0/FzqRPI2rJt9GrwRsp9TgwYj5OejiCkvC4tJLy7nClhB8249
PbkmTP2j+kXMCp8H5b/FW8bLg+4+agl/oAcwWvP03b43nkIMqt/YUBtUEkIzPi2C
ZHjckic+OpeoVNLeDUkpUhbu4hCH2YeENm6JTaw3fME=
`protect END_PROTECTED
