`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC2o2Sg9PmNHP81pXPokLqxEjUaQSLEvJYi3OVtz4K6+
ZteP3cg7wMbvidN2RYA0L74klrxtFs4Vfdj51RiOg45dCnk7jTG6LmmTJ2Ly0sh7
P2cCUubmTBQzfMziaOOw7LvGGwsknZL141uaHFky5oyzyTW9ueqFLBbfId7TgJJp
aa2E8TYsbuc6SLYGb7lOYTH3qZJ+K1FGzW6D8WdHc4m8fhVCzYOrH8Vl6eQqLyS0
`protect END_PROTECTED
