`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKA2OMuHQHS6Sn0Rt3qiNPoWM6mlexX4DBv+cmVKNknC
7fPccIhTSSpCpm+IzuHNgXsPYIf3SLl3UB9maKx6IBcuahq89H/t6dEQeGM3YDew
dlDb2qh4qjWa4YYGXRN78jqEBbOtH8mOurhNIkTIjsREgDd2Zi6pDJLC+cLAm6VB
/5U7Iy1H1UZ7ayVgCOEvrmpH4CLymuS8/vx86KlVCcXtgjAvZ/eNcnSQkjcCB4Ta
DA+p7DHAsDJucDq7yd2w2Z3vGsM0kiJQIN9c2iljPBy0ic+3GmwFy3c8O45Lj8pE
YoN8PVBwK9fOwJEeXbZLOOQDs/2Jm89/9ut7wI8IjtnwavKcKO9EO6+GJ1AVQGcY
fsT1hjFPVG0SyF4JCDY5VqQPQcl4ydtKqHEPO0eWQWHqC7Neo6EieRkCW2TH7VxT
8K5We8tOb+jEJbuEwbYgeLzOq680CUXIrxMzymJTUsVOtvq0lqgQossTlKVI5VcE
JcPvyOffq75XWRTroCz7iTZlSzHa9qkQbmyrDRnwJLW32gz6wp2f9PITAVT6fe3w
vEA9zxCKhHObv6/wN+7iDQ==
`protect END_PROTECTED
