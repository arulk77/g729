`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNjeTbtJrKsCq3EosTHeA5xMg+5sA8kOB0DTveA1ttVg
pYhBWlovDjZGyY2nNJhM+qjuQFlvmJ7O9IBkicdT/sdh6ajeaFxAitLOCur4WxLS
v5QcdncGSDOTJb7caKCa6Y5sqAjnZqqpL41t1hJrRC9dsZcr54qZ/vAE1oPU4sfk
g8714WC5FypsBvkNQX/K7WyX8BAqm7PxgBsh5/d0ZZE4JTh+Iaai1GgOeGd8LybV
8ulM2SpRsQSpSFt0m9c/oCwo1vUiYbvJr2+OPLXDVrsU7LjymbizGxcIbg0C1CZ0
NtoCIXDbV2ApWm2TiYsxnNmEgoxn1LQdcAPAwi0BacrIBmAhv1kGFCJgZR+Z67dn
ouv5k8sxGZg0cJezYkQoDQ==
`protect END_PROTECTED
