`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePYHUDVaQ6i7Sn1LNqspcvZnvWMIt4YS8ZCosxcNNKnc
v7Fuqq9AcjCzzFlEDsuEC0hu7kikpv1n0DAwXQzyAJwcCH9IqptxQsz8YM3PkMnm
mLegXVuStRDL7LwqcuXgvXFySSg5LmDwgg7YkeBNGCQfUl8JxNKENj8B7v1OTUTr
rSSpgJfF9n0ecDKNi4K2131VmzheGziMc9giA8MYbAWVAQuxYyjIJJhHFiDGccZf
HwYVbXbb6qAlvBcI9tU3TqT9FTpj2SW681bPsB1m3JcjfrkpamKzOVELcR10c98x
KzyJKN/IcH53+xA3/czkkg==
`protect END_PROTECTED
