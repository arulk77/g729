`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL0O0FgWq1Zrzf1gulofLxLPux+UU4hfT0MLYfNnvdQN
5MLoR2i9m3c1Yj3oF8jOjvYjxOXiXSu+H37j9TjUwCgq+O/BQ2h6MaKVoNjoe8UE
UhLSrlvhEN0GOiIZDEeA17/TX5l+s9I5Us9J7wUv6zSso6Gt5DGbRBY5s+lRhDml
5ilhFu61QTUGIx3bYPFzOLk3SvG7I/BeplpRMjgVtipe1KcfqJVk8wpAcCECfMnU
bML1EO1vKcI8wyC6CQ5XgIa3izC2J8eHGzxtUCXl+WixonGLsuL6C55ERAbJSyKi
uWUo/54N2iKXWH9fWZKF5JnHK0bKL/ySaMItayyucetC1NtRYV1YtTnj+ojXWTec
xwMb03IV48sJWRyZZlofrhpZxKrq6OGg6yd5pMFfncBnGkkRQyEB4ueRoERveFR7
Bh8/ZgqdLz/09unL0t8JB++HyAPqZChRpwSBp8bzzvmP3SufGNmW3jTJB3nBS2en
Q58bAeZVsDTux38qU3fRUZbaB9DVX0aZHRWKcIGSn/V5Y2W8PIX0dRz3nS6yU5W5
PD6kb0D3VfeYfGLac20cOA==
`protect END_PROTECTED
