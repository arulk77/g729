`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+QGUATRrOeEBM4ICu33oxYMraEvP6hVYChU0uCD1Gcn
2AFFzXil+3tDsrK8WmRkb5IQkd9mWstcqL1vvJVS+FHVcSSpQt2x4MO10Wo42uDP
TT01g1lCZbUGMsThwH3PmyKP8wCSEZqmyHAh+Qx8nN2s0bwyiLVJLpQxfx/JmoZm
2fnumq5Q3Gu5qAUvizsXP78i0WDyLwBBbTalNHmMh1s=
`protect END_PROTECTED
