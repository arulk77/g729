`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abD4Id8uSOw0bMPEDWQjU3QHQM9UQglHBvyyFRs68erR
DLdi01oQ1E9BmEkhKOBAW0vt5vhfYbxytLjWg9wZTZ9/OmxrGRr1ygbm3AlNna96
4cCIy2G9ywfxkHvivRI90+CJtVHY07aTaN8Wmz5Df6XjUpONSDm97f+FFn6LP3et
To83eP6u6k8Lms4wGktTkEfQMRce54VN/qPw6FK3bqj7pYId5u6y5sBuliq66cuJ
FCN1htHKNOn5CjgmgBvm+xZsOWG0IRtCKYYKz4oyt5HaTmeA0hOeK0U6F4klDP7S
mFjj4poErE0tN4z5T3kHJIxJTXApjqGn7rDr53a5kJmhZCozbWaxf1fTgh086FDO
NqoPtZPgDk0bEj2AWaVCT2L9OEmv9w25xRWEVZEhw/Le3dQCdtAZpoKEVxcHm0Eg
8KNsu1s9gqzyTKDhPxFSBY8k314C8IM7v3dqrtX6Xxtw9fTCZkEdruhg/pnKGK64
H95J1Tq0I0/gLhszCwNMCaaxzoRReHCJO12JKRqd/2ZqK4eJm702a9X8oM5x1nZE
TiRXmPeXFP2E7VNF0ezMNomy2feM9lDQu8DEmwSDTGwsK68zMbBZegpZ6jHxrZhe
ifRcnwTREWOr+2Q97PHe3l5uRiafA3duGhNvYfkVbyB+blE4I6eipWOqYsvLC5kp
/CHHf9V0RUc/X0FVtoS6SBcr9qJQCaFDowlx9XrAvAtX1KRsjjifIcKAiIDwq81j
sl4/tiQ9RNZ1kloGoD5jrzkG7U0+KXFXMk0UIjKn1nyg/SvIBe2g/dYYPmKZZP9R
sq+1MuE6dva57QuQDFZqrUxSs+FlihqO9lIqvG5EWk1x61duu17sjSQ5XrRr/BPJ
Xkwtbf2yzHhhj2FZar92EnsPog9IvngfqFwmS5zUGECuE24+PEurTIouu13Xh6Y0
jcl25t36iuzgnNBWF5LOCKl5BqXy2EYz8yB3RQ3Q+Ksmmsg7c0omsBeKUOxhlKMR
3TQiyaINaxz8ia/cBlfELrBJgpj5pfZPS4WYDru27atcNEtzhlHVceJ6iGtS+6ZL
JE2mBU9yNKDZjDtGZwukbFYTkTbgy8BRX0rgZOomYQE4Um9psdmxaDQTxk1TZ3jD
ZKFqkpokPIGyH/jgzZwiGCAZqcyKoWPPmjjOsCXHc53Q3CFZ+GOFrSOYL8qQbfSB
AiSXvq5uE3uistQfkMz8g3jZwG+HC5Y2rOl6dv6ox0bbC9gxn22dOGaAk2p6Hpyt
GR9U3bqLRUuJyVo5GC/Wsy+ovIxcRTD3jFbbdIba5OOGrItWG5akhKEKeMGDIV2S
1+W8Nvijalcs3AWdX4lyCXbzSRWZssQKU1CTl4F3nUP72ptWP9AIEjEu64V8ijlu
KS6G7f8olyj6M+aZ/qQ/fm74hcyo2LamJQwCT4EpA341Homoaca0X3gjHjKLLZMA
fpShsGwHLcpKcr+to3kj+vy7rqJize0BjOyLqf6DpokGaDAiwnmaHpHsoxOLbw9d
jGGzLHxH4xHwcyine/BdaWRE2h8IMvKztGpehUHQHyLzjPC5vIHtB7XahWmjIiiI
XdP9BT8dhIXKg8M3Sg1OpE3pC1yPrAVxfg742I79+1eh3Qvu5KFjyxxVnP+O1zyt
Ry6FJM5wykE2Dc8Oz12/jx4DpAoOLrRVSKd5VP61ATPee0a7zgDy1PM6uYn8Yptz
LQzLregfLNVyA1XiBW6Jl7VC7oClaBUKmhVpubyK7WJNdTlGyGoZK7vtl0Qcmm4I
UbPQf7wTgVMPQxFIv+NrpAp5t+7UaZJ9gzf2VZ+HkMgQOLbbcdrggTkw7/JBg5gJ
uNK1cyZX9BmicW6QvVhd14ZTL8WevdWVyjRiZ/SpTTOq+VF82pEbFpdlhn4K2tNZ
7InkCJWqvVMNIHUPpsQUQih337nkusUaMRVlCqNIaKnopSkiyzWynYcM9BuraHaM
4KTDh6Xo9LQMTsGz/3SpU5zgloYuAFrPufN6VXLYeqNYVDrzWTTvwjxjQ73MI4DK
9ejLTa5Jb6p92rhLHKIbrQamnFyFNYvJfbvbCzr7WGR7a4Im3KKybNyftjzPu6tn
bMR6+2PXItW3FBa0K0MH0crSMT24X5rSFsIvD5tNwWdAyXcXUMKdAw7Ug44Qv7Ha
IZ9yX5e6JyuabKniE6dWGLrs6H0Zj8uaU2AdWYK9La2dLpjVR8t91Pi86bZAd7go
vqhqEyciKvBGS8EmbhwfUCEhYaVgvWVsCZBcIp08T784ZsRQhoOZ5MgDcAzRyrwx
61KlS5T6Lqw3O0W3i8T6zGJYi/JTMj/2Qi/20+dvql8s4+jRGcKXOjYkJ399JkW0
GO4NgS579gZK0YNLyRD6phwtELtbGreseTeFv1LLifVery159UXgLXlX6a5OS+xL
7/8r2ywkBi5zezBhosuwLzYaSObqEP/bZxThsp+AUE215ivtWFJDgOplkl9P5ZQq
rUf1KUv8B2k8qBEbYujg5GbuBnbuPbHoIgMYzp+U2/dIqbbEtao0a8P0r1oTK8Ke
2rR7+buv6y/xaXefq4oCQcW2O+L4uNjufsFJlntPoDxGK15nB6My+cC4pBfVXRej
OyBGUrDTxH2zQkpusrW8X4JrauXP7sAGwaHN2rzLxY2JuGIxg2GVmUdmNrYfLxwo
pKU1yKdTAEHYxkBLMjzCygHuEM+fyU7UCQ+6ojEaaLY9OPPkevZc12KQg86/wflA
lDaiLBSzOev/Zoyf1FR4fKZq+NoSBQMeflV83IxdXBPVWf4Fo1QYUUkYip725SRf
xLHkWc4g7O5ii8BR1ULKfhRUCmXPJHwK7tigsZW8IlS+QrUeOQC26A0JEFU6J75y
OKhZCfizbgvg7+Tk+cdR93Y/qWBCpQV9SOJCA3439IbpQJxy0LUWXGOTZvHXOo60
usbHeRSj7v7BivzieqVoptIgUFXEaKaaNLK4H42XSIJS3xsDbJM0glXRBPvkJ1eg
lqVwUA1NawaEfe9uesoD5FhaYNIcpKoAoJFnK08xwaMtnCZAxHGD0VcbI8vE0Asn
vJRHEHy1anpLXL3yldkQhJ6EwVl9JHGx+IBq5UIfzzk3wBPuouvjb2XDjz3/mq9B
I0h5uEbMSy+V9LSWl6WM2GA1P3f+T9dnhDJI2O4tYsXCGnlWNMI5bcnBOGmLRSdb
4UeJZHYNvs8C6GfMqbqq5pZ+nU75ppbI/UWL09T40BOUU8Hh8kNtieVlScUhCDX3
Q4LtDb0jtsp6GI5k3iNfITo9w69gf2EZ/fpyjW2iotHkesAy33x2p/vAAsn6GJ5Q
M3zA6wSGAUldlZGP5uj5PSa+VD7fEtoOpUSPXyjBgCsz5xFm8jF/dlbUou5vs++K
VKOnjk0uqfveZ+E5HrHa3iEm3rwycvn1Z81Vcb9zfqT27dSzcHhfUP7oMncs1rgR
pcxU55O16DJadyxp+VoCz6aDQCrWIR0QohXByUo4/NH4rhzMxi3ULPNPVu28qPP+
FZSEPHKkeMCF1qlLBycBOC6q6hXR9KshPxDxT9cNk0jsOerAutkO024CH4gEn4Sr
d2z61Xx8wpS6otuEwS9EdNZZ74ZCK23jGFa6N8kWl1avoqQdWDjQfMNDZdJI4rvH
LHMMRckYNQnhLs40n+oXD6Fh4EFRvYoQzHSsxAOSWeQRsHTH3RdcsVcor24ftnPD
z2HCPrzDBMxqo03C0iEcrUPHmBdx/OUM21MYRpnyYDq9dN+Suo38l6MYqqIusYVW
OhPHuG/lQlZVRfKQSUrycbXW/4OJ+L1YsARDoXChfcPCFBxPw7kj/ZIRhxS70vKh
Hsb8YS0KbKO9TflDNeXnv0qycRn70x58R5femVSVSiBvdYwf9bzPZxKhnSYT5N4v
mrtb9enccjOp2SlNIoLrpR8UPzCVk7Rxgjoi5Qn8ywMbNWKbS2eEErDgV02syXe7
uMsPJMKSRo0b8Zol23QJWVMO0dxo/0nTNmrlpbFhuihSW/zJZstpDt4r+XI5gTdq
3s/K7Rn51VaHQ09+5h2e/M3XoiPvfBDNYa+4BJ1E4XaYWqr96sECauJ88avROUF9
HZLf0ETzUlA2i/ZPTPqCVg2W3ePwj/q2/3q0Pk3oTu8STM+8d8RdEezt0mo+rjUZ
h1Iqs4EZfInw0/303OS7OjOCGvcoN0OsQenGuDBzrEZJHc6j5v9og+wqvcwX2VJZ
+hYTTUNC1QkkQSXg9Nu2UnzVPgGbFI5jeBcTfO7ZEbbhXHEhA42FkWzEM+2VsZaZ
Af4VdokVaCfTh+LNnHCTxjpirmot3HSZ9ZpbrfRz6v6oXky+mvocBdCITkxN6Kxy
N7yMhvjzqjVUXPhz+2xIw09oe38gJ6nK68JZD6lbLBPINLzdoK9kCsshvZypaAA3
Y0nTjGWDYEC1u2vkzw9pjtXo6+EXM42WpY/KZlIT3rpEhMLYCwOjgPpS4BQDskTk
yobFxPuIhbWEco+yj4xG38MPas08h6/jYIz/JP2lrjz2jz+fxDw2ZyJBXtbQ3b/Y
gO5o8kVnI13YmJuzuFDnyZuJFrvjR9giC7VKVrVk2KWXz57wgqYpbl52YqTDbbT6
sja08Jtn58K0MA6J17d1pjH0aCiX1V9HdxvGL1yvWp31pkWTYJ4MG1aHX3iDTchD
6qkC7AGjLUOV7uNEPm1mReM7ICJGWwA6rcat4eLs+V2K0vTb+rEJZ8yNRfTclG+3
BK+mNpwxyqS+o+vUeNv38qx/h/hX3fsKL+43/sC0OV/VLIHQ6CTnxOWaRoFzWtJU
6pHYI0aWBHh6oY2905Lw1e3gGD+P59hdR23vOHLWkZq1kf3SO8xj9XMeLpxdBJ7I
FrFYIHYFecZKaf1FjD69fti6v48a0vQw3qwIxBrAUS5u0hZ0qjiK66JAlfm7kxJq
K7WkA+4FlTrPAuPGGos0KDYIQUxGUqjHlE63FkSZVMmFwQBBf/rv2fz/llCYrXFn
r1zcJMAKj98UnzhNN2byUdls9ZcW3WXVhMq5+PiAIidxZPaBSelashyYQooNWvd0
gM8jt8EUfmQZdhzOaEiORBDy8JC9pzmo2eqfvqkf4QvM6ducaE/V2e4SCCFvcqVz
l6Ba5gjouvq8Uq5Evfu4ucDBEIRAO/P3TkkVyLi8TAZ0IKHwpTB9/jV8OB1Kkpbp
AtcIFzSoDt2tyMJbbnFszDK0zziz31JNxQrCT1BqU0xTAIAW3nCf8otg5zKpvPDl
Fx/2IazyVV06dAsxNuffyCGNNI7TvEj7jFBZoVY1tWLaCo9deMBpdbsDVbWa9rR8
WjVG4n+D85lUpMESKTLsXd21mqXcfCG4UGATkqel7wc3zIHx69S/KQK/urvKPuJO
VoHps2tUXMb0YpS7qVn7BRycITpGaO0w238hsdxCO+hY25Fark6HA3ghHHPg31TT
lkxZ0IeaI63ZOoZEOo+S0UJgtb815HdsBFe3xcAg1Bw0Ln8pcZvzBL0GYYphrxWI
jKsdpg6WgPQMd60cEIgzPxwFHgoP6hphTqYxz7dh4yHOlKRQP25MMfl7WGzgETUH
hqKS9cjR77KdYARTWg1rt8zA/4b2cPUvjbtvQhPfhWUt2XqAJtt5F3QuUtWJGg59
2Z8xCRBRev0TBjT4fXcx1Upszsp8earFE/K2rOKYXhu6Ed/VjL8vDsZx8Z6FdgF6
uV0fhPhu5O3I6OkqoyfWuisctmKOh0S8IVI36e9KLE9HjVCVggKMkxYj8dK0lJl8
PvpU4A73JcxNS3wAPdexpdJYz5vHRDH7/E5B0/9IGLEZYr1/bHIqHH9yMBfK8aSZ
96T/M/NZUlnHk3eps/TeNHtZ15E0wMstZ1wPqgrGh0nRGlx2c7OeozLoqwtyHvkl
NC4b016drc6ZRqKIK6r4ahVaSU33GZx5GC2Yzb55WrGxLSGHD0bnbm1DByclU414
r9+aNPmvpu2B0hNC2Hn3QJNl8jqx2nEliNwauzeL4igs70g5OOGon0m7NVS3dmnL
UbK4cQaalbSfoTqnXbpL6j/BjqSzKjpvEk2YvuZWsRlNHGEZ1y83dYL2BzFSjHN9
L8ZHOGe3i4i6OFangxSWpqrqgaq6q5UD+4CMp41zYgDioqIOITCRfoPoK9g+vFRl
BVO/bCJ6cupCvzOVwRWlZm1fmv5mFxaWUUZXYW7j4NNNGRK6KVSojnwsr/ffGO9g
NHe2n3bjWEiZZ0e3yUoXbaiFAEdE1deGQ8aUVSlSkVl7lmlzR4qjWucxJXIkWmfY
D7Tc/EgDSM60PM28xy+r3eW3dZMcuApuQHotdZKUaA0l1pmkE4jUsxIesNWzgVom
8c4p14KtjlkKoAIlKFHxB9pqb6Vxk/l8lvNp5cdRHkskMacpP9LPtPy4Afvkjzjp
JGPCjRRILhK8AhKLx404lOSYjwGgK3ETEU+jU9IjSTagNt0dmkj/B/m4aunfq50v
cA3iaRDUV1yTCbaX45Am71f9M9+aefJty/5zVkHpr9l0cpXasd+JqSmq1i5GdcZT
7syojRDSsRtcHgrymLIUVKEiO81slgqOmlThdzY6XJvE0cW+NCPGj2Z2eV4ZwglJ
yJ37nkPzN0ps4Bvh/mOi4ZEFowGaciDVcsxABHxmtpBBzGpP+M9BrrraaIPin6cM
+ZvL3ksLJ6ALw/qtUZAbtJj2o/Qrh6IblXl/GVv3zfygbVK1sbVeh0VcAOXdL2+9
QWTMDnw3Pbd9CmdvjnPvA1EJblmmL/+2E6tZNeVm3dx2o+TH0uDDKqeCMKkrUm4F
7B2YW5T9xzTuqLYEIKTwaVF/q1lqeN7mLir7iLRRX4E+JMak34YofDSGOc/MHMVo
IO+zbba7BytBEBNYzU6pMlBG7BZeVoqUZ8uKfHTrKaDklmVhI9UOxnE4QBGhrHsS
8npPWs8/MEtvx9SpmSd3oq2nEbztJ9cz4mcxyzv4Qa1fLvzhoUkfk4WoPKcJskCK
Zh1Mln1X5OcPGxdcoz+OdIBZmlCxM7oZD87HS5F9gDRBESz3cQ6/2LmQb8lj4+h/
L3TgNBGBE8nX25Px3j4dZ1Ea9/ksxxjplihJOL53uHPNBZk8QCW79hF2bmGy5aBC
G6sk3lnCPIfh+hr8EpfOQWl+FDmqEJAJwgmy+HevOCjKq+s8uQpCMyAbPc9p1QCU
U/sSMjD/pEnLWg8Ym8P9i6jVWJPoySjW9p2kbx6zYqStY3JG5QSkAxQETh319shg
YOvKj9dx/FUrld2N7s6kSdPor0e31amr2hsotd1v6QM+8V5HlF4zhYFigBvG0nnN
z8LcDz/6vRQIHEAENg7LwnP8jVwbV9Ad+KdxPLn/HOg5UxA9Ey47D2sTakpjADXE
jQbxuGzumOU7h0VruOI7bA5SYS/dO0BI+r6bt1gDv/w3hshwhC8mcywpkOmaWsSZ
UNqxzUqM1QNKP10+HOqfoe2bpgPG6b/QAfFZO8ySov9411XQNWWSzW7kswmc0JtC
lFWnhQnjjDSFntZOkHOnWQQpFll8oIVVjhQpT6GQT7TulfAaN3ua6Zr2xb45pD5m
t8bi1RCotKzcbZ61nnuxuyFyTS3MkQ8y1JUWzBZcLNwnFhbPjZt11h8APlKbLORk
HRfP0XEkwbDKwo+9qmPGT/VAdftUle1HbZn0PAkmuD7nA/e56HuBypxEZQMQjhMc
u3M6ZJTL8wZJnAzQ1xtpnqqD202kBoqpipw4If41154DGGY6z/nvZ7EaK8Z58OaM
c/DZO4HEHPm2k3RNW4OVxWszJ97WiLdhxwbjjCemHL2mk7AkPGzEfGHLIDjmtmHU
+nfPQ7Gl/qpUDC/BVZ0pKnUZ0HzfusnlXE2WV68Y0Zser7dKoeDQfp2wllqugK4o
E8krG7Dx86Rw7SYlQnUuquegLVzH7k1KH/gyeQwsEUNmFSNeMfnkgOie4jAOglt1
A81sJR/owD6vN3FcNG9MYUirxzav7nsr5hapzlOoex1pTkV2ozoJNVE9QOCQP8Cp
4ZheQD4MbTiYOKQfF3oOAHO9hK7bhG/VO4TDbs7BRqaaximpdVqkkR4hou+nv7pq
/qb8vBhrWuNLI0Q7hJnn4/RIGp63i7LbSnOO2b7LlUuqaAcv0qxZ9U4yGrFtevGb
mvQotfpIpZnASweDzbBy8ZKp7/p/BGeko4k9AXVVn3zGBgZGY3DqIicmBfjX2vik
PPEZJ/EcXPuex++tCAy4Kxfin8cW+E2uqwnytslZWDAN5vNb2xNS0tsOFg05CekY
sdBhX0yksr6p+anRSAAcap8Bc0AfG4BsU9US4QGmYO3hPn/VHmv8xi0/VziVuWJB
ukhmCsgnJZ6n+3b7AHFNSghAui8+753Cv9TtbaZiuAemnqCpD2saedTVDSqlsntZ
qL24U2RpQGXVWK6vaFWlG3DngUhur885NBwHm+XuU0vU6aK1OuXZU6IKZNkXnmjN
b32WwFTiFSRPTKvDpOmjyfbQmMJ9ZU059kveWiWjEMZTEUFxaMAl8lBW8iXatUQF
20PW9yEJU4RIPX8feitUTI1CpoTMytbzxY/M64+t3XujYBETbc+RztC0g98OcuaZ
3zt33deVFtnl40vc51pFGiKJs7B97yWsEmHdyac5gQUKYM99s7tRNrBw9ElZbepU
U8tLurobE+yBJK2Bv+LLhy0zQprW5iQOGAX8/1XCHAk1f2/R5SyMoBMOFbNIMk+m
f2FMuCY3h821dpO6GayAuniwHvLxmKmwxRVdJI5rKPKhYaR7k2+I0Mah/Z4c6zu5
6lZyc7z5x6Xdpcw4+IXHmvE8uf1Rtx5pYrLCXC+zqNbSAFaxBEtCStolzpH8YJgI
nk1wYI6wGxekLJGmYTXwWjAwfKrkKejaQxk56K6LP1Y+4V8QX/8ym/Hgg0DYHfyz
Hym+UbXShIDqMlwQD+lXL506U+8IgLFnko7YULXfLm3jNZTTmHtbkGgFfmq+3EFo
mK6bCmZgAOIuRZysk5j4I82jpKw8uvd3hMGjfABlwqICrYd4C8WEPQFIQyPkFCU1
5zcgHs/MGO75/DQ9Lu9NpL6Dh4QF2u2gwvolsONdTuYLBfxjAf2tHenLrBk1v8hy
QafzbJ1vkmH1fzyoZEGlpYOQ3bGIVqDUuhX761hs7D0e9MJbHyP0UVZ5vaLa25Xd
riayCl1Rk+vk/nZnwocK+rFpxjUyBPvK3/NvqImQP13ztHl7VFFgnAb4JO1sNfC5
Na/lAWzQllBD3OLbqR3t139s/PaSIGawOB0+0kXLsKEX+in25j+edrwI/L+qyhVD
MzYB6W5Agp25UnSeVG5wNAsyfsFNaRQ8ZYkCljwgr6o5XxUBRuQZHZcKpsNnkNr2
Ed6XDFYFlL3Eo3fgiKgx/q+P+zkSVinTGCzGvUI/x17kU+aBrkKoQYU5khsE2irv
jhn36c0SQImKpboRqsUI5EP5Ja+D0A5lXN0Mc0XsBckTImyb1T4W5YEOaZBxUPtp
+a1xzPl72OaPb4ENR5oXXvpepGAo9rVOHC+vZSpn4cnL46eDf8jMeVEazXaXAL2e
CqPFo5BlT2TPzZnmbtMWvHTV5rcxkQ9zo+2WYFs7hP9u6UKuaVGNwMHCFFLIVJb3
wYKFhlYVtWGiV1MXhBK4x2IhAAf858+qCtbhIySXqKdbRlWAbCVWaGWnOB0WpwJb
+IKbVGfnrrIukhwuz4bLEeXj5bNfac23LIefcoYCWz2UGoAII/RHVLB6t2lSr9pg
e11FicFvDn0AuG/FzTsQOP+jkRm4fR0FRAp3StrXVAL4Zn7o7nTY1zQq3J7WCSbt
MrLxohwa1/oRn0noYP6k1vYNNa6B76DFMORcHHmRh0zC5CunwQVXcW+u2YHFPlcu
HSGq1l9LTON1xCed1vmruHAdTXBDbhh+olHyEbBM2j4mYlpagxkSrtgFRxlXG80N
qYRM1DKfRqo3tMno7ZQmhI8Pe5KasR6rJYR2GpxGl/xzxmpFFySl23mdyADTPgpU
Ocks3IyHw5ISqdcpYa6yJu3iS3PNLXTKrSszauWuwbKnF88tfzcov/+R9P4fnGz2
UcFRqd7xi3CfzSy1uVC7j9jtsSuwtTkciC+pxUMHJxLDeSFUzjePhbdmW84oat7n
M1SKaOl0/ya3CK704l00+JFmpSWdVl3GvawED8pRYMNRzGHcUtzMfWFJX4dswRzl
`protect END_PROTECTED
