`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAL/pG3SF5svpCWAyjQMp9L+c5ZJHmbYcQ+SNJd7RVQa
Am396eVurY/+SWUDibVJ41Q6+M+XA5FTEVfNq9GMznaiAat5Wa6IX8UQcK+7yWCe
fTFib/lrTw2aBposyt4/GNCIVS5KiW+xsK22sJjOcbHfwi451ZMo9Pd5uXlG9fFy
qvTmz7RG7oorseT4kmbruRpKynqWzXZXWOKwn7NlgwmrZxQEn4LfoyoDNkLzkVfJ
XUXQd6h+RgLMFUtPTnR8DkKwFtQeqdtN/bZWdjUqQ3SG3cKVOHbKZXhzfQMks8WZ
eg2bK058dlxFJUqBf7y7wQ==
`protect END_PROTECTED
