`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49cX5HTRFwlHvlXd87AHsZNb5pnwNHyreyR7s7NJ8bNv
xiwjX5Zs1MkQ6uYqCXxdf0py6ds/oxRvpw9dxd5BGF77fycyDKv7+1/+sc7cu+/2
/hDUOSO12vF485+3tVQdbbEKcMHETuyaJH1yW3QZbMuf75BF4fBD7UuEd5dA9y6c
IivP/oKefncROTUKOJ5yJw+D4hJBJx+UOy4I1nYr/hX2lhJFQM5RN4ACPicWRvLW
thf+4jcvZ5CbAX8WLdxqcZlx/+S3SIAD9WIo7pkr+YY9biY7vAKDH6TJ1ZgzVE5c
zA7HQhAov5A1A21t1eTWkwH6yjBPcfBGH0ZkHSy2fuwpHJK6K+RBp/0D36g+qAoQ
EKwRAyd0o8hNPWwm3ZAkHA==
`protect END_PROTECTED
