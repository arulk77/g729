`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePLsHht4gVwNfQyBxy52/Ak0UhIlZnEGQ34zedtW7mBR
FhaI8CM7kZKdiatKWsXVcy5iwiEzhWN3lIfij9Ui3p3W8sRwyJjPdgNzVrnA8Sg9
0ficLD4rlywKwJnBFoUbW+5C/YEPJkTRv2N/16/uFZJdwbjWW+ABh2Sd8DRHWh0D
L3sixi5iCsmF8oUy7n3DZDM3LJIgc1dj7JU089gGuDFvkLmWs4Xuzq/SIgtitRba
KIomXNSugnhWqMoQiOM6CRKazf+zDlpIsmAoSao/7zLd3N2BIOXg1GUCvxTD6EsK
J6DmjpMIGyY0lp/7+KFuZf+r/dDK21XCO4iS0AwpJ+zWW2uOrFMuSWRXGfaDds6f
ja8O6d4OJB+ELvpPjoeaMvn5KZqs+CxsAfOMj5t46hHGzNf77BGczQDBe8UqX51O
88LkF7nwQ5XQzroVTXq+zwi1xO0Haas4H93aTO+sfKtOjylU5oxP/i/w5VJ/8iJx
Xc3MI4s87tqnOwZcEbJxfD/tiZDEpuBSk7dAMjzuKNiB6TOtJhXh7JFbQmB6gdJB
`protect END_PROTECTED
