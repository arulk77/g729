`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
v5FiHTHsrFLJopN/RMgg7yTF9nIGDQoPenzdTZ3mrZPLPbtBbDQqvS8g0ZwKqoER
W4KtaUA6UNvGheoYzRXkd/SHBPVdi09HYGtJ9KrScKPrnDlDXI2cibEmKwhcHACa
8FIibsA9opVyJjSNCJd029RefSH+0GpXYrZZhuXr7klu35Hs6yxWV/XASHZ4uOaW
l2DLA9RSHay1SpZVtpC5Nr7PxFCOWFj7ZVAv8s5gjWiOPXIjb6CiIXRfMyxvNuvR
QR9km1AMpPpG++7TjmgjqgdhR/qUZZPJe4TYdvIBpaLP3AAJ3sKKScFJuJv8D9k+
Zds+ZtceoCRT4ne4EumJaREn1JFDXf2JyiSQ/HYTv6kkufeZJjYUaswie+5ltD7f
L6c5V/z9EXft4E0Qvuzel+YSJnrEkfNOTO6YWC5Ef61Aa09jJIzcVWruUWCd3vwL
YNl8kWtiFmvGDjHMdpWMYRDRjNtau9Xgkyg4N9LfTPNV1ax4bex6j2Os4LCysbxW
49YirnXXUpv5NM/eLV7nxbzgJCN9Q4GlN1dxx19Gf3TK2GUknzfWppDbiMxji1a2
7yhtTSjt5XpOIVDEZI4+uYjQvkPCk4DreF2eHfp2PdGG9PnF2CRDlSPM8iVSIfbS
DOb7H2fkvLwm62W+45o6u5mS9euiUNYaysjFZi9YuooIVL6+mweKa48qDCRLWZDa
`protect END_PROTECTED
