`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
oUBIC3HaU3aM4AbVDC0rGbwru9xocAFjAqQjJyz2/N1sV4JUJXqGb034DV4QS3y4
wR1U0tdmPLA0oSlmh8bflq/2vcKRO3IttFmZvLMUcEqgXerSwUooTXSM9uoJ5srW
dwDYtmtaHDHctQyEnvFPalnf4vqBDVNaQLHuob73qeA23djWNjUMCE6JN8dP9Vi7
huDGh/3VgUaTlm8mqRNjTxchhgP9c8plhxmDcZ4go8CZLaQu/5VvRUx6FllYeEFC
CI2pUCexmOhr6k62YlZJS0KLraa8rMHJMPMyZ+otZKmS4BcYnUsa/enyY7ZuMEbv
+ovvrvPN7CdwIVP6T7kc61cxh2diJfSi0UxHB5I+pJ/EsGnyB8hh0NdJ0sbwjEhg
PwlVF+0hBhkwjL5Fsw+vxJq6xinczxSu2wU7t1EobsA=
`protect END_PROTECTED
