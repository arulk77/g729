`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49vLVpsJZIBsU7UbIdLoKxf8iHs0NA5DhKe91coNSVH0
/Kbx9cEdprR7LRw2AfYNey2qa2d20p/MuMeY1+EViWMhaEz9bRPUz0rzkRGWC7e7
JIF0qhDv9/QamOGIb6+36fxT6NBAPEMy4UfTrKJbwteEq94Q/bFSO//NHzIU/X3l
CVV1ICLd272nHMryz5dwB3Fitb+vGRJl4l/xgona1/U=
`protect END_PROTECTED
