`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yKJYz6kU6tJlOvHARWajoams3V6+Jv2idz86NMSVxVF
6rT9KkpS+Fku+6LmIcE+LZwFO/ChA76lWOduVXBdSFttlUZwSQMRxVkBjL4GMySH
uVWVWXruwqmi8U04EjZ3LGpDkJG2hWIrm9x9g6Ka56WfKBVWku51WMI767NSmdNy
jsUls1Z1FyvlBCz985BwAC+Ql2A0iGEMP2SBLpvRpxUOf55ataOpvSWDmOtYQRC+
+cMuaihDzvR7SzGX+o+Vrmnj69tboT9YWbXIHGgNSn3mC8LDq8wkFQqWjEiGUIkN
OnZGcMTLnJWE86j85/yxxImBw7gjaAYHv9fIMdcqQ6TOsZBcTVLU8yoEsr9Mwkkv
Rge0xymYcVMastWc3V+DfQ==
`protect END_PROTECTED
