`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN2yGGfdJcMRAFzHfnpWgPtjDo7Ia/5OrBKfFaYb4wBRW
c5D7mR7nGuMkj18Z5YiFLtd7U3rDXvAnhWoqcVUd2IMvVE9ntvTSJtSHOraArhWM
2whNbckhBqNfQwb8/YTm5O//tsFZsoD6EkD6rpaKQfbBPcJbc7jhly28Gd5Xqteh
EYrCrbQDoXX362pGKvpJWuqMWr61oTKIYjKiGslRBnL094cCbT+KfU0haZ/bKd6e
ffC/2XC3iSsoF/nFbfwS5segihRDaT2MbjX4iX2BeiMImG4Qb9NV3HAeh6h8zlbq
sjf0FMLRFnI4psh0r5PlsVCn1lnR8MLQYhlAbOekcXkInU0veBGg2fEtDR7jsp2k
EKXLeHRDR3zxycaRBWXv39wvyaOrnLLsspB0DGm7Xk2X0KYXwX7CaXyhOTHteRKr
Y/I9E2M1H0wE1Tx/XbzqkacZzT1ZwOSB/PGlToNhEQUSk0EQNGUn6htkKOW/X+Vm
AUCMDf3LRwYnG6HHEGJI2FHFqmeNHqBAL3jBaPjzNPD7QUu81Z2i2ytv3hcsp2VF
/P/FgddZm2PQcZ/qaqQUT4mUzK88zRXVcUJ1rpK6QegsWpsFTlxAbB8AwBBFX5OF
zw7+3gojlms6eM09Fop6dHal73AnFgzqF6WtzhQhkSuS4eumWZ9GSL7PtKgHq8oT
0Xv9sIs1VUc1uZb8x5DyQcBVkT+nZmYduS3giJUkboBED+Xazg2XKIFSXcECuE8w
AcCIQ6BB09TJ/hOGy0Kt7yLwjUbdFH1SukJxBeI/SnZ+tUCSvY0kePqRXwTlxlTz
m8Hi9ICwFU9tg3Pl5RYeESsXJtRpIe4wxnZ3c7PQj+lSMq9U9Od97kByPTqxgQkF
g5qWreF5vB5Y1GgWQQfNpBikErvsVI3a1eF1JU0jGME=
`protect END_PROTECTED
