`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDRzk4JCpeEOAHCcDVOj/jjVy1UfGWyjkVY/YNUZNuCz
YoAtuyPynRZ1ekaWx7PoT9icv9I0p9+Imj/eyefDKVERz65QUhATt1bTMNk2/Jig
LIQOpBMrGKl2zd3fN9Pn9VsS5wKVmfPYPXRkwNLFP3w64sz0hEt/DjQOCanwIM51
BKk9Pc6/j2NhckLuDwGrpRmz1N5qf5Gu/jy9h37WAT1M6ZTNU/siTypJxY9B+kjg
Zp97qgNSXlYZ8BvWcRaIJQNQ2xAjH0/CqVwqhyHxVGpeorWmGsL4X1L+r/wlCyox
9cWOu5nTNuCFVxpuewpgZ3QPt6HLWGGJtRmrOkKYMKfENxxLwaW+vFJ11kd9SR46
Hg7VOuoFqI9lrcK0ag5HMb0+/kphSRvGHNHgcZ+xrvE=
`protect END_PROTECTED
